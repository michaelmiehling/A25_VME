-- z126_01_ru_cyclonev_m25p128.vhd

-- Generated using ACDS version 14.0 209 at 2014.11.19.13:38:25

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity z126_01_ru_cyclonev_m25p128 is
	port (
		read_param  : in  std_logic                     := '0';             --  read_param.read_param
		param       : in  std_logic_vector(2 downto 0)  := (others => '0'); --       param.param
		reconfig    : in  std_logic                     := '0';             --    reconfig.reconfig
		reset_timer : in  std_logic                     := '0';             -- reset_timer.reset_timer
		clock       : in  std_logic                     := '0';             --       clock.clk
		reset       : in  std_logic                     := '0';             --       reset.reset
		busy        : out std_logic;                                        --        busy.busy
		data_out    : out std_logic_vector(23 downto 0);                    --    data_out.data_out
		write_param : in  std_logic                     := '0';             -- write_param.write_param
		data_in     : in  std_logic_vector(23 downto 0) := (others => '0')  --     data_in.data_in
	);
end entity z126_01_ru_cyclonev_m25p128;

architecture rtl of z126_01_ru_cyclonev_m25p128 is
	component z126_01_ru_cyclonev_m25p128_remote_update_0 is
		port (
			read_param  : in  std_logic                     := 'X';             -- read_param
			param       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- param
			reconfig    : in  std_logic                     := 'X';             -- reconfig
			reset_timer : in  std_logic                     := 'X';             -- reset_timer
			clock       : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			busy        : out std_logic;                                        -- busy
			data_out    : out std_logic_vector(23 downto 0);                    -- data_out
			write_param : in  std_logic                     := 'X';             -- write_param
			data_in     : in  std_logic_vector(23 downto 0) := (others => 'X')  -- data_in
		);
	end component z126_01_ru_cyclonev_m25p128_remote_update_0;

begin

	remote_update_0 : component z126_01_ru_cyclonev_m25p128_remote_update_0
		port map (
			read_param  => read_param,  --  read_param.read_param
			param       => param,       --       param.param
			reconfig    => reconfig,    --    reconfig.reconfig
			reset_timer => reset_timer, -- reset_timer.reset_timer
			clock       => clock,       --       clock.clk
			reset       => reset,       --       reset.reset
			busy        => busy,        --        busy.busy
			data_out    => data_out,    --    data_out.data_out
			write_param => write_param, -- write_param.write_param
			data_in     => data_in      --     data_in.data_in
		);

end architecture rtl; -- of z126_01_ru_cyclonev_m25p128
