-- megafunction wizard: %ALTGX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: alt_c3gxb 

-- ============================================================
-- File Name: Hard_IP_x4_serdes.vhd
-- Megafunction Name(s):
-- 			alt_c3gxb
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 15.1.0 Build 185 10/21/2015 SJ Standard Edition
-- ************************************************************


--Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus Prime License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


--alt_c3gxb CBX_AUTO_BLACKBOX="ALL" device_family="Cyclone IV GX" effective_data_rate="2500 Mbps" elec_idle_infer_enable="false" enable_0ppm="false" equalization_setting=5 equalizer_dcgain_setting=1 gxb_powerdown_width=1 hip_enable="true" loopback_mode="none" number_of_channels=4 number_of_quads=1 operation_mode="duplex" pll_bandwidth_type="auto" pll_control_width=1 pll_divide_by="2" pll_inclk_period=10000 pll_multiply_by="25" pll_pfd_fb_mode="internal" preemphasis_ctrl_1stposttap_setting=1 protocol="pcie" receiver_termination="OCT_100_OHMS" reconfig_calibration="true" reconfig_dprio_mode=0 reconfig_pll_control_width=1 rx_8b_10b_mode="normal" rx_align_pattern="0101111100" rx_align_pattern_length=10 rx_allow_align_polarity_inversion="false" rx_allow_pipe_polarity_inversion="true" rx_bitslip_enable="false" rx_byte_ordering_mode="none" rx_cdrctrl_enable="true" rx_channel_bonding="x4" rx_channel_width=8 rx_common_mode="0.82v" rx_datapath_protocol="pipe" rx_deskew_pattern="0" rx_digitalreset_port_width=1 rx_dwidth_factor=1 rx_enable_bit_reversal="false" rx_enable_lock_to_data_sig="false" rx_enable_lock_to_refclk_sig="false" rx_enable_second_order_loop="false" rx_enable_self_test_mode="false" rx_force_signal_detect="false" rx_loop_1_digital_filter=8 rx_ppmselect=8 rx_rate_match_fifo_mode="normal" rx_rate_match_pattern1="11010000111010000011" rx_rate_match_pattern2="00101111000101111100" rx_rate_match_pattern_size=20 rx_run_length=40 rx_run_length_enable="true" rx_signal_detect_loss_threshold=3 rx_signal_detect_threshold=4 rx_signal_detect_valid_threshold=14 rx_use_align_state_machine="true" rx_use_clkout="false" rx_use_coreclk="false" rx_use_deskew_fifo="false" rx_use_double_data_mode="false" rx_use_external_termination="false" rx_use_pipe8b10binvpolarity="true" rx_word_aligner_num_byte=1 starting_channel_number=0 top_module_name="Hard_IP_x4_serdes" transmitter_termination="OCT_100_OHMS" tx_8b_10b_mode="normal" tx_allow_polarity_inversion="false" tx_bitslip_enable="false" tx_channel_bonding="x4" tx_channel_width=8 tx_clkout_width=4 tx_common_mode="0.65v" tx_digitalreset_port_width=1 tx_dwidth_factor=1 tx_enable_bit_reversal="false" tx_enable_self_test_mode="false" tx_slew_rate="low" tx_transmit_protocol="pipe" tx_use_coreclk="false" tx_use_double_data_mode="false" tx_use_external_termination="false" use_calibration_block="true" vod_ctrl_setting=4 cal_blk_clk coreclkout fixedclk gxb_powerdown hip_tx_clkout pipe8b10binvpolarity pipedatavalid pipeelecidle pipephydonestatus pipestatus pll_areset pll_inclk pll_locked powerdn reconfig_clk reconfig_fromgxb reconfig_togxb rx_analogreset rx_ctrldetect rx_datain rx_dataout rx_digitalreset rx_elecidleinfersel rx_freqlocked rx_patterndetect rx_syncstatus tx_ctrlenable tx_datain tx_dataout tx_detectrxloop tx_digitalreset tx_forcedispcompliance tx_forceelecidle intended_device_family="Cyclone IV GX"
--VERSION_BEGIN 15.1 cbx_alt_c3gxb 2015:10:21:18:09:22:SJ cbx_altclkbuf 2015:10:21:18:09:22:SJ cbx_altiobuf_bidir 2015:10:21:18:09:22:SJ cbx_altiobuf_in 2015:10:21:18:09:22:SJ cbx_altiobuf_out 2015:10:21:18:09:22:SJ cbx_altpll 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_counter 2015:10:21:18:09:23:SJ cbx_lpm_decode 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_stingray 2015:10:21:18:09:22:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_stratixiii 2015:10:21:18:09:23:SJ cbx_stratixv 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY cycloneiv_hssi;
 USE cycloneiv_hssi.all;

--synthesis_resources = altpll 1 cycloneiv_hssi_calibration_block 1 cycloneiv_hssi_cmu 1 cycloneiv_hssi_rx_pcs 4 cycloneiv_hssi_rx_pma 4 cycloneiv_hssi_tx_pcs 4 cycloneiv_hssi_tx_pma 4 reg 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Hard_IP_x4_serdes_alt_c3gxb_41f8 IS 
	 GENERIC 
	 (
		starting_channel_number	:	NATURAL := 0
	 );
	 PORT 
	 ( 
		 cal_blk_clk	:	IN  STD_LOGIC := '0';
		 coreclkout	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 fixedclk	:	IN  STD_LOGIC := '0';
		 gxb_powerdown	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0');
		 hip_tx_clkout	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 pipe8b10binvpolarity	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
		 pipedatavalid	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 pipeelecidle	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 pipephydonestatus	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 pipestatus	:	OUT  STD_LOGIC_VECTOR (11 DOWNTO 0);
		 pll_areset	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0');
		 pll_inclk	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 pll_locked	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 powerdn	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 reconfig_clk	:	IN  STD_LOGIC := '0';
		 reconfig_fromgxb	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 reconfig_togxb	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => 'Z');
		 rx_analogreset	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0');
		 rx_ctrldetect	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 rx_datain	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => 'Z');
		 rx_dataout	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 rx_digitalreset	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0');
		 rx_elecidleinfersel	:	IN  STD_LOGIC_VECTOR (11 DOWNTO 0) := (OTHERS => '0');
		 rx_freqlocked	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 rx_patterndetect	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 rx_syncstatus	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 tx_ctrlenable	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
		 tx_datain	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
		 tx_dataout	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 tx_detectrxloop	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
		 tx_digitalreset	:	IN  STD_LOGIC_VECTOR (0 DOWNTO 0) := (OTHERS => '0');
		 tx_forcedispcompliance	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
		 tx_forceelecidle	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END Hard_IP_x4_serdes_alt_c3gxb_41f8;

 ARCHITECTURE RTL OF Hard_IP_x4_serdes_alt_c3gxb_41f8 IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "suppress_da_rule_internal=c104";

	 SIGNAL  wire_pll0_areset	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_pll_areset_range50w51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pll0_clk	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_pll0_fref	:	STD_LOGIC;
	 SIGNAL  wire_pll0_icdrclk	:	STD_LOGIC;
	 SIGNAL  wire_pll0_inclk	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_pll0_locked	:	STD_LOGIC;
	 SIGNAL  wire_cal_blk0_nonusertocmu	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_adet	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_coreclkout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_dpriodisableout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_dprioout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_fixedclk	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_quadresetout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_rdalign	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_refclkout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_rxanalogreset	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxanalogresetout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxcrupowerdown	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxctrl	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxdatain	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxdatavalid	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxdigitalreset	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxdigitalresetout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxibpowerdown	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxpcsdprioin	:	STD_LOGIC_VECTOR (1599 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxpcsdprioout	:	STD_LOGIC_VECTOR (1599 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxphfifox4byteselout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_rxphfifox4rdenableout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_rxphfifox4wrclkout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_rxphfifox4wrenableout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_rxpmadprioin	:	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxpmadprioout	:	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxpowerdown	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_rxrunningdisp	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_syncstatus	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txanalogresetout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txctrl	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdatain	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdetectrxpowerdown	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdigitalreset	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdigitalresetout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txdividerpowerdown	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txobpowerdown	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txpcsdprioin	:	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txpcsdprioout	:	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txphfifox4byteselout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_txphfifox4rdclkout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_txphfifox4rdenableout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_txphfifox4wrenableout	:	STD_LOGIC;
	 SIGNAL  wire_cent_unit0_txpmadprioin	:	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  wire_cent_unit0_txpmadprioout	:	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  wire_receive_pcs0_cdrctrlearlyeios	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_cdrctrllocktorefclkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_coreclkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_dprioout	:	STD_LOGIC_VECTOR (399 DOWNTO 0);
	 SIGNAL  wire_receive_pcs0_hipdataout	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_receive_pcs0_hipdatavalid	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_hipelecidle	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_hipelecidleinfersel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_receive_pcs0_hipphydonestatus	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_hipstatus	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_receive_pcs0_parallelfdbk	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_receive_pcs0_phfifordenableout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_phfiforesetout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_phfifowrdisableout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs0_revparallelfdbkdata	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_receive_pcs0_xgmdatain	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_receive_pcs1_cdrctrlearlyeios	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs1_cdrctrllocktorefclkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs1_coreclkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs1_dprioout	:	STD_LOGIC_VECTOR (399 DOWNTO 0);
	 SIGNAL  wire_receive_pcs1_hipdataout	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_receive_pcs1_hipdatavalid	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs1_hipelecidle	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs1_hipelecidleinfersel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_receive_pcs1_hipphydonestatus	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs1_hipstatus	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_receive_pcs1_parallelfdbk	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_receive_pcs1_phfifordenableout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs1_phfiforesetout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs1_phfifowrdisableout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs1_revparallelfdbkdata	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_receive_pcs1_xgmdatain	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_receive_pcs2_cdrctrlearlyeios	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs2_cdrctrllocktorefclkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs2_coreclkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs2_dprioout	:	STD_LOGIC_VECTOR (399 DOWNTO 0);
	 SIGNAL  wire_receive_pcs2_hipdataout	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_receive_pcs2_hipdatavalid	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs2_hipelecidle	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs2_hipelecidleinfersel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_receive_pcs2_hipphydonestatus	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs2_hipstatus	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_receive_pcs2_parallelfdbk	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_receive_pcs2_phfifordenableout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs2_phfiforesetout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs2_phfifowrdisableout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs2_revparallelfdbkdata	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_receive_pcs2_xgmdatain	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_receive_pcs3_cdrctrlearlyeios	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs3_cdrctrllocktorefclkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs3_coreclkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs3_dprioout	:	STD_LOGIC_VECTOR (399 DOWNTO 0);
	 SIGNAL  wire_receive_pcs3_hipdataout	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_receive_pcs3_hipdatavalid	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs3_hipelecidle	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs3_hipelecidleinfersel	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_receive_pcs3_hipphydonestatus	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs3_hipstatus	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_receive_pcs3_parallelfdbk	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_receive_pcs3_phfifordenableout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs3_phfiforesetout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs3_phfifowrdisableout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pcs3_revparallelfdbkdata	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_receive_pcs3_xgmdatain	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_receive_pma0_w_lg_freqlocked613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_receive_pma0_analogtestbus	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_receive_pma0_clockout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma0_diagnosticlpbkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma0_dprioout	:	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  wire_receive_pma0_freqlocked	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma0_locktodata	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_reconfig_togxb_busy514w601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_receive_pma0_locktorefout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma0_recoverdataout	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_receive_pma0_reverselpbkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma0_signaldetect	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma0_testbussel	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_receive_pma1_w_lg_freqlocked681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_receive_pma1_analogtestbus	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_receive_pma1_clockout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma1_diagnosticlpbkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma1_dprioout	:	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  wire_receive_pma1_freqlocked	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma1_locktodata	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_reconfig_togxb_busy514w677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_receive_pma1_locktorefout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma1_recoverdataout	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_receive_pma1_reverselpbkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma1_signaldetect	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma1_testbussel	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_receive_pma2_w_lg_freqlocked748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_receive_pma2_analogtestbus	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_receive_pma2_clockout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma2_diagnosticlpbkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma2_dprioout	:	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  wire_receive_pma2_freqlocked	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma2_locktodata	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_reconfig_togxb_busy514w744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_receive_pma2_locktorefout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma2_recoverdataout	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_receive_pma2_reverselpbkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma2_signaldetect	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma2_testbussel	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_receive_pma3_w_lg_freqlocked815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_receive_pma3_analogtestbus	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_receive_pma3_clockout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma3_diagnosticlpbkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma3_dprioout	:	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  wire_receive_pma3_freqlocked	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma3_locktodata	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_reconfig_togxb_busy514w811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_receive_pma3_locktorefout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma3_recoverdataout	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_receive_pma3_reverselpbkout	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma3_signaldetect	:	STD_LOGIC;
	 SIGNAL  wire_receive_pma3_testbussel	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_coreclkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs0_ctrlenable	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_datainfull	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_dataout	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_dispval	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_dprioout	:	STD_LOGIC_VECTOR (149 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_forcedisp	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_forceelecidleout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs0_grayelecidleinferselout	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_hipdatain	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_phfiforddisableout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs0_phfiforesetout	:	STD_LOGIC;
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs0_phfifowrenableout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs0_pipeenrevparallellpbkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs0_pipepowerdownout	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_pipepowerstateout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs0_txdetectrx	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs1_coreclkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs1_ctrlenable	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_datainfull	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_dataout	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_dispval	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_dprioout	:	STD_LOGIC_VECTOR (149 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_forcedisp	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_forceelecidleout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs1_grayelecidleinferselout	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_hipdatain	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_phfiforddisableout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs1_phfiforesetout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs1_phfifowrenableout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs1_pipeenrevparallellpbkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs1_pipepowerdownout	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_pipepowerstateout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs1_txdetectrx	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs2_coreclkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs2_ctrlenable	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_datainfull	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_dataout	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_dispval	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_dprioout	:	STD_LOGIC_VECTOR (149 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_forcedisp	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_forceelecidleout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs2_grayelecidleinferselout	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_hipdatain	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_phfiforddisableout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs2_phfiforesetout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs2_phfifowrenableout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs2_pipeenrevparallellpbkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs2_pipepowerdownout	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_pipepowerstateout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs2_txdetectrx	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs3_coreclkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs3_ctrlenable	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_datainfull	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_dataout	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_dispval	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_dprioout	:	STD_LOGIC_VECTOR (149 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_forcedisp	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_forceelecidleout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs3_grayelecidleinferselout	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_hipdatain	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_phfiforddisableout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs3_phfiforesetout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs3_phfifowrenableout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs3_pipeenrevparallellpbkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pcs3_pipepowerdownout	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_pipepowerstateout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_transmit_pcs3_txdetectrx	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_clockout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_datain	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_dataout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_dprioout	:	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  wire_transmit_pma0_rxdetectvalidout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_rxfoundout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma0_seriallpbkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma1_clockout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma1_datain	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pma1_dataout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma1_dprioout	:	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  wire_transmit_pma1_rxdetectvalidout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma1_rxfoundout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma1_seriallpbkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma2_clockout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma2_datain	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pma2_dataout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma2_dprioout	:	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  wire_transmit_pma2_rxdetectvalidout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma2_rxfoundout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma2_seriallpbkout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma3_clockout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma3_datain	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_transmit_pma3_dataout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma3_dprioout	:	STD_LOGIC_VECTOR (299 DOWNTO 0);
	 SIGNAL  wire_transmit_pma3_rxdetectvalidout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma3_rxfoundout	:	STD_LOGIC;
	 SIGNAL  wire_transmit_pma3_seriallpbkout	:	STD_LOGIC;
	 SIGNAL	 fixedclk_div	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 reconfig_togxb_busy_reg	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_w_lg_w_lg_w_lg_fixedclk_sel57w58w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_fixedclk_sel57w64w65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_fixedclk_sel57w69w70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_fixedclk_sel57w74w75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_fixedclk_sel53w54w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_fixedclk_sel57w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_fixedclk_sel57w64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_fixedclk_sel57w69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_fixedclk_sel57w74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_fixedclk_sel53w54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_reconfig_togxb_busy514w515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_fixedclk_sel57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_fixedclk_enable52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_fixedclk_sel53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reconfig_togxb_busy514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_analogreset_range513w612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_fixedclk_sel57w58w59w60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_fixedclk_sel57w64w65w66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_fixedclk_sel57w69w70w71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_fixedclk_sel57w74w75w76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  cal_blk_powerdown	:	STD_LOGIC;
	 SIGNAL  cent_unit_quadresetout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  cent_unit_rxcrupowerdn :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  cent_unit_rxibpowerdn :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  cent_unit_rxpcsdprioin :	STD_LOGIC_VECTOR (1599 DOWNTO 0);
	 SIGNAL  cent_unit_rxpcsdprioout :	STD_LOGIC_VECTOR (1599 DOWNTO 0);
	 SIGNAL  cent_unit_rxpmadprioin :	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  cent_unit_rxpmadprioout :	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  cent_unit_tx_dprioin :	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  cent_unit_txdetectrxpowerdn :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  cent_unit_txdividerpowerdown :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  cent_unit_txdprioout :	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  cent_unit_txobpowerdn :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  cent_unit_txpmadprioin :	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  cent_unit_txpmadprioout :	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  coreclkout_wire :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  fixedclk_div_in :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  fixedclk_enable :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  fixedclk_fast	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  fixedclk_sel :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  fixedclk_to_cmu :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_pipeenrevparallellpbkfromtx :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_rx_coreclkout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_rx_phfifordenableout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_rx_phfiforesetout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_rx_phfifowrdisableout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_rx_phfifoxnbytesel :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_rx_phfifoxnrdenable :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_rx_phfifoxnwrclk :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_rx_phfifoxnwrenable :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_rxcoreclk :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_rxphfifordenable :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_rxphfiforeset :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_rxphfifox4byteselout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_rxphfifox4rdenableout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_rxphfifox4wrclkout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_rxphfifox4wrenableout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_tx_coreclkout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_tx_phfiforddisableout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_tx_phfiforesetout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_tx_phfifowrenableout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_tx_phfifoxnbytesel :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_tx_phfifoxnrdclk :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_tx_phfifoxnrdenable :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_tx_phfifoxnwrenable :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  int_txcoreclk :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_txphfiforddisable :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_txphfiforeset :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_txphfifowrenable :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_txphfifox4byteselout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_txphfifox4rdclkout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_txphfifox4rdenableout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  int_txphfifox4wrenableout :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  nonusertocmu_out :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  pipedatavalid_out :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  pipeelecidle_out :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  pll_powerdown	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  reconfig_togxb_busy :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  reconfig_togxb_disable :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  reconfig_togxb_in :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  reconfig_togxb_load :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  refclk_pma :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rx_analogreset_in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_analogreset_out :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_deserclock_in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_digitalreset_in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_digitalreset_out :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_enapatternalign	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_locktodata	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_locktorefclk_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_out_wire :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  rx_pcs_rxfound_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rx_pcsdprioin_wire :	STD_LOGIC_VECTOR (1599 DOWNTO 0);
	 SIGNAL  rx_pcsdprioout :	STD_LOGIC_VECTOR (1599 DOWNTO 0);
	 SIGNAL  rx_phfifordenable	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_phfiforeset	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_phfifowrdisable	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_pll_pfdrefclkout_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_pma_analogtestbus :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  rx_pma_clockout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_pma_recoverdataout_wire :	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  rx_pmadprioin_wire :	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  rx_pmadprioout :	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  rx_powerdown	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_powerdown_in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_prbscidenable	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_reverselpbkout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_revparallelfdbkdata :	STD_LOGIC_VECTOR (79 DOWNTO 0);
	 SIGNAL  rx_rmfiforeset	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rx_signaldetect_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  rxphfifowrdisable :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  tx_analogreset_out :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_clkout_int_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_datain_wire :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  tx_dataout_pcs_to_pma :	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  tx_diagnosticlpbkin :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_digitalreset_in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_digitalreset_out :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_dprioin_wire :	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  tx_invpolarity	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_localrefclk :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_pcs_forceelecidleout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_phfiforeset	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_pipepowerdownout :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  tx_pipepowerstateout :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  tx_pma_fastrefclk0in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_pma_refclk0in :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_pma_refclk0inpulse :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_pmadprioin_wire :	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  tx_pmadprioout :	STD_LOGIC_VECTOR (1199 DOWNTO 0);
	 SIGNAL  tx_revparallellpbken	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_rxdetectvalidout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_rxfoundout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_serialloopbackout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_txdprioout :	STD_LOGIC_VECTOR (599 DOWNTO 0);
	 SIGNAL  txdataout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  txdetectrxout :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_cent_unit_dpriodisableout1w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_fixedclk_fast_range56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_fixedclk_fast_range63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_fixedclk_fast_range68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_fixedclk_fast_range73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_analogreset_range513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  altpll
	 GENERIC 
	 (
		bandwidth_type	:	STRING := "AUTO";
		clk0_divide_by	:	NATURAL := 1;
		clk0_multiply_by	:	NATURAL := 1;
		clk1_divide_by	:	NATURAL := 1;
		clk1_multiply_by	:	NATURAL := 1;
		clk2_divide_by	:	NATURAL := 1;
		clk2_duty_cycle	:	NATURAL := 50;
		clk2_multiply_by	:	NATURAL := 1;
		DPA_DIVIDE_BY	:	NATURAL := 1;
		DPA_MULTIPLY_BY	:	NATURAL := 0;
		inclk0_input_frequency	:	NATURAL := 0;
		operation_mode	:	STRING := "normal";
		INTENDED_DEVICE_FAMILY	:	STRING := "Cyclone IV GX"
	 );
	 PORT
	 ( 
		areset	:	IN  STD_LOGIC := '0';
		clk	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0);
		fref	:	OUT  STD_LOGIC;
		icdrclk	:	OUT  STD_LOGIC;
		inclk	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		locked	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneiv_hssi_calibration_block
	 GENERIC 
	 (
		cont_cal_mode	:	STRING := "false";
		enable_rx_cal_tw	:	STRING := "false";
		enable_tx_cal_tw	:	STRING := "false";
		rtest	:	STRING := "false";
		rx_cal_wt_value	:	NATURAL := 0;
		send_rx_cal_status	:	STRING := "false";
		tx_cal_wt_value	:	NATURAL := 1;
		lpm_type	:	STRING := "cycloneiv_hssi_calibration_block"
	 );
	 PORT
	 ( 
		calibrationstatus	:	OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		clk	:	IN STD_LOGIC := '0';
		nonusertocmu	:	OUT STD_LOGIC;
		powerdn	:	IN STD_LOGIC := '0';
		testctrl	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneiv_hssi_cmu
	 GENERIC 
	 (
		auto_spd_deassert_ph_fifo_rst_count	:	NATURAL := 0;
		auto_spd_phystatus_notify_count	:	NATURAL := 0;
		coreclk_out_gated_by_quad_reset	:	STRING := "false";
		devaddr	:	NATURAL := 1;
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		in_xaui_mode	:	STRING := "false";
		portaddr	:	NATURAL := 1;
		rx0_channel_bonding	:	STRING := "none";
		rx0_clk1_mux_select	:	STRING := "recovered clock";
		rx0_clk2_mux_select	:	STRING := "recovered clock";
		rx0_clk_pd_enable	:	STRING := "false";
		rx0_logical_to_physical_mapping	:	NATURAL := 0;
		rx0_ph_fifo_reg_mode	:	STRING := "false";
		rx0_ph_fifo_reset_enable	:	STRING := "false";
		rx0_ph_fifo_user_ctrl_enable	:	STRING := "false";
		rx0_rd_clk_mux_select	:	STRING := "int clock";
		rx0_recovered_clk_mux_select	:	STRING := "recovered clock";
		rx0_reset_clock_output_during_digital_reset	:	STRING := "false";
		rx0_use_double_data_mode	:	STRING := "false";
		rx1_logical_to_physical_mapping	:	NATURAL := 1;
		rx2_logical_to_physical_mapping	:	NATURAL := 2;
		rx3_logical_to_physical_mapping	:	NATURAL := 3;
		rx_xaui_sm_backward_compatible_enable	:	STRING := "false";
		select_refclk_dig	:	STRING := "false";
		tx0_channel_bonding	:	STRING := "none";
		tx0_clk_pd_enable	:	STRING := "false";
		tx0_logical_to_physical_mapping	:	NATURAL := 0;
		tx0_ph_fifo_reset_enable	:	STRING := "false";
		tx0_ph_fifo_user_ctrl_enable	:	STRING := "false";
		tx0_rd_clk_mux_select	:	STRING := "local";
		tx0_reset_clock_output_during_digital_reset	:	STRING := "false";
		tx0_use_double_data_mode	:	STRING := "false";
		tx0_wr_clk_mux_select	:	STRING := "int_clk";
		tx1_logical_to_physical_mapping	:	NATURAL := 1;
		tx2_logical_to_physical_mapping	:	NATURAL := 2;
		tx3_logical_to_physical_mapping	:	NATURAL := 3;
		tx_xaui_sm_backward_compatible_enable	:	STRING := "false";
		use_coreclk_out_post_divider	:	STRING := "false";
		use_deskew_fifo	:	STRING := "false";
		lpm_type	:	STRING := "cycloneiv_hssi_cmu"
	 );
	 PORT
	 ( 
		adet	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		alignstatus	:	OUT STD_LOGIC;
		coreclkout	:	OUT STD_LOGIC;
		digitaltestout	:	OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		dpclk	:	IN STD_LOGIC := '0';
		dpriodisable	:	IN STD_LOGIC := '1';
		dpriodisableout	:	OUT STD_LOGIC;
		dprioin	:	IN STD_LOGIC := '0';
		dprioload	:	IN STD_LOGIC := '0';
		dpriooe	:	OUT STD_LOGIC;
		dprioout	:	OUT STD_LOGIC;
		enabledeskew	:	OUT STD_LOGIC;
		fiforesetrd	:	OUT STD_LOGIC;
		fixedclk	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		nonuserfromcal	:	IN STD_LOGIC := '0';
		pmacramtest	:	IN STD_LOGIC := '0';
		quadreset	:	IN STD_LOGIC := '0';
		quadresetout	:	OUT STD_LOGIC;
		rdalign	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rdenablesync	:	IN STD_LOGIC := '1';
		recovclk	:	IN STD_LOGIC := '0';
		refclkdig	:	IN STD_LOGIC := '0';
		refclkout	:	OUT STD_LOGIC;
		rxanalogreset	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxanalogresetout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxcoreclk	:	IN STD_LOGIC := '0';
		rxcrupowerdown	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxctrl	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxctrlout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxdatain	:	IN STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
		rxdataout	:	OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		rxdatavalid	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxdigitalreset	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxdigitalresetout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxibpowerdown	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		rxpcsdprioin	:	IN STD_LOGIC_VECTOR(1599 DOWNTO 0) := (OTHERS => '0');
		rxpcsdprioout	:	OUT STD_LOGIC_VECTOR(1599 DOWNTO 0);
		rxphfifordenable	:	IN STD_LOGIC := '1';
		rxphfiforeset	:	IN STD_LOGIC := '0';
		rxphfifowrdisable	:	IN STD_LOGIC := '0';
		rxphfifox4byteselout	:	OUT STD_LOGIC;
		rxphfifox4rdenableout	:	OUT STD_LOGIC;
		rxphfifox4wrclkout	:	OUT STD_LOGIC;
		rxphfifox4wrenableout	:	OUT STD_LOGIC;
		rxpmadprioin	:	IN STD_LOGIC_VECTOR(1199 DOWNTO 0) := (OTHERS => '0');
		rxpmadprioout	:	OUT STD_LOGIC_VECTOR(1199 DOWNTO 0);
		rxpowerdown	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		rxrunningdisp	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		scanclk	:	IN STD_LOGIC := '0';
		scanmode	:	IN STD_LOGIC := '0';
		scanshift	:	IN STD_LOGIC := '0';
		syncstatus	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		testin	:	IN STD_LOGIC_VECTOR(1999 DOWNTO 0) := (OTHERS => '0');
		testout	:	OUT STD_LOGIC_VECTOR(2399 DOWNTO 0);
		txanalogresetout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txclk	:	IN STD_LOGIC := '0';
		txcoreclk	:	IN STD_LOGIC := '0';
		txctrl	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		txctrlout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txdatain	:	IN STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
		txdataout	:	OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		txdetectrxpowerdown	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txdigitalreset	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		txdigitalresetout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txdividerpowerdown	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txobpowerdown	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		txpcsdprioin	:	IN STD_LOGIC_VECTOR(599 DOWNTO 0) := (OTHERS => '0');
		txpcsdprioout	:	OUT STD_LOGIC_VECTOR(599 DOWNTO 0);
		txphfiforddisable	:	IN STD_LOGIC := '0';
		txphfiforeset	:	IN STD_LOGIC := '0';
		txphfifowrenable	:	IN STD_LOGIC := '0';
		txphfifox4byteselout	:	OUT STD_LOGIC;
		txphfifox4rdclkout	:	OUT STD_LOGIC;
		txphfifox4rdenableout	:	OUT STD_LOGIC;
		txphfifox4wrenableout	:	OUT STD_LOGIC;
		txpmadprioin	:	IN STD_LOGIC_VECTOR(1199 DOWNTO 0) := (OTHERS => '0');
		txpmadprioout	:	OUT STD_LOGIC_VECTOR(1199 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneiv_hssi_rx_pcs
	 GENERIC 
	 (
		align_ordered_set_based	:	STRING := "false";
		align_pattern	:	STRING := "UNUSED";
		align_pattern_length	:	NATURAL := 7;
		align_to_deskew_pattern_pos_disp_only	:	STRING := "false";
		allow_align_polarity_inversion	:	STRING := "false";
		allow_pipe_polarity_inversion	:	STRING := "false";
		auto_spd_deassert_ph_fifo_rst_count	:	NATURAL := 0;
		auto_spd_phystatus_notify_count	:	NATURAL := 0;
		bit_slip_enable	:	STRING := "false";
		byte_order_back_compat_enable	:	STRING := "false";
		byte_order_invalid_code_or_run_disp_error	:	STRING := "false";
		byte_order_mode	:	STRING := "none";
		byte_order_pad_pattern	:	STRING := "UNUSED";
		byte_order_pattern	:	STRING := "UNUSED";
		byte_order_pld_ctrl_enable	:	STRING := "false";
		cdrctrl_bypass_ppm_detector_cycle	:	NATURAL := 0;
		cdrctrl_cid_mode_enable	:	STRING := "false";
		cdrctrl_enable	:	STRING := "false";
		cdrctrl_mask_cycle	:	NATURAL := 0;
		cdrctrl_min_lock_to_ref_cycle	:	NATURAL := 0;
		cdrctrl_rxvalid_mask	:	STRING := "false";
		channel_bonding	:	STRING := "none";
		channel_number	:	NATURAL := 0;
		channel_width	:	NATURAL := 8;
		clk1_mux_select	:	STRING := "recovered clock";
		clk2_mux_select	:	STRING := "recovered clock";
		core_clock_0ppm	:	STRING := "false";
		datapath_low_latency_mode	:	STRING := "false";
		datapath_protocol	:	STRING := "basic";
		dec_8b_10b_compatibility_mode	:	STRING := "false";
		dec_8b_10b_mode	:	STRING := "none";
		deskew_pattern	:	STRING := "UNUSED";
		disable_auto_idle_insertion	:	STRING := "false";
		disable_running_disp_in_word_align	:	STRING := "false";
		disallow_kchar_after_pattern_ordered_set	:	STRING := "false";
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		elec_idle_eios_detect_priority_over_eidle_disable	:	STRING := "false";
		elec_idle_gen1_sigdet_enable	:	STRING := "false";
		elec_idle_infer_enable	:	STRING := "false";
		elec_idle_num_com_detect	:	NATURAL := 0;
		enable_bit_reversal	:	STRING := "false";
		enable_self_test_mode	:	STRING := "false";
		error_from_wa_or_8b_10b_select	:	STRING := "false";
		force_signal_detect_dig	:	STRING := "false";
		hip_enable	:	STRING := "false";
		infiniband_invalid_code	:	NATURAL := 0;
		insert_pad_on_underflow	:	STRING := "false";
		logical_channel_address	:	NATURAL := 0;
		num_align_code_groups_in_ordered_set	:	NATURAL := 0;
		num_align_cons_good_data	:	NATURAL := 1;
		num_align_cons_pat	:	NATURAL := 1;
		num_align_loss_sync_error	:	NATURAL := 1;
		ph_fifo_low_latency_enable	:	STRING := "false";
		ph_fifo_reg_mode	:	STRING := "false";
		ph_fifo_reset_enable	:	STRING := "false";
		ph_fifo_user_ctrl_enable	:	STRING := "false";
		phystatus_delay	:	NATURAL := 0;
		phystatus_reset_toggle	:	STRING := "false";
		pipe_auto_speed_nego_enable	:	STRING := "false";
		prbs_all_one_detect	:	STRING := "false";
		prbs_cid_pattern	:	STRING := "false";
		prbs_cid_pattern_length	:	NATURAL := 0;
		protocol_hint	:	STRING := "basic";
		rate_match_back_to_back	:	STRING := "false";
		rate_match_delete_threshold	:	NATURAL := 0;
		rate_match_empty_threshold	:	NATURAL := 0;
		rate_match_fifo_mode	:	STRING := "false";
		rate_match_full_threshold	:	NATURAL := 0;
		rate_match_insert_threshold	:	NATURAL := 0;
		rate_match_ordered_set_based	:	STRING := "false";
		rate_match_pattern1	:	STRING := "UNUSED";
		rate_match_pattern2	:	STRING := "UNUSED";
		rate_match_pattern_size	:	NATURAL := 10;
		rate_match_pipe_enable	:	STRING := "false";
		rate_match_reset_enable	:	STRING := "false";
		rate_match_skip_set_based	:	STRING := "false";
		rate_match_start_threshold	:	NATURAL := 0;
		rd_clk_mux_select	:	STRING := "int clock";
		recovered_clk_mux_select	:	STRING := "recovered clock";
		reset_clock_output_during_digital_reset	:	STRING := "false";
		run_length	:	NATURAL := 4;
		run_length_enable	:	STRING := "false";
		rx_detect_bypass	:	STRING := "false";
		rx_phfifo_wait_cnt	:	NATURAL := 0;
		rxstatus_error_report_mode	:	NATURAL := 0;
		self_test_mode	:	STRING := "prbs7";
		test_bus_sel	:	NATURAL := 0;
		use_alignment_state_machine	:	STRING := "false";
		use_deskew_fifo	:	STRING := "false";
		use_double_data_mode	:	STRING := "false";
		use_parallel_loopback	:	STRING := "false";
		lpm_type	:	STRING := "cycloneiv_hssi_rx_pcs"
	 );
	 PORT
	 ( 
		a1a2size	:	IN STD_LOGIC := '0';
		a1a2sizeout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		a1detect	:	OUT STD_LOGIC;
		a2detect	:	OUT STD_LOGIC;
		adetectdeskew	:	OUT STD_LOGIC;
		alignstatus	:	IN STD_LOGIC := '0';
		alignstatussync	:	IN STD_LOGIC := '0';
		alignstatussyncout	:	OUT STD_LOGIC;
		bistdone	:	OUT STD_LOGIC;
		bisterr	:	OUT STD_LOGIC;
		bitslip	:	IN STD_LOGIC := '0';
		bitslipboundaryselectout	:	OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
		byteorderalignstatus	:	OUT STD_LOGIC;
		cdrctrlearlyeios	:	OUT STD_LOGIC;
		cdrctrllocktorefcl	:	IN STD_LOGIC := '0';
		cdrctrllocktorefclkout	:	OUT STD_LOGIC;
		clkout	:	OUT STD_LOGIC;
		coreclk	:	IN STD_LOGIC := '0';
		coreclkout	:	OUT STD_LOGIC;
		ctrldetect	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		datain	:	IN STD_LOGIC_VECTOR(9 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT STD_LOGIC_VECTOR(19 DOWNTO 0);
		dataoutfull	:	OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		digitalreset	:	IN STD_LOGIC := '0';
		disperr	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		dpriodisable	:	IN STD_LOGIC := '1';
		dprioin	:	IN STD_LOGIC_VECTOR(399 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(399 DOWNTO 0);
		elecidleinfersel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		enabledeskew	:	IN STD_LOGIC := '0';
		enabyteord	:	IN STD_LOGIC := '0';
		enapatternalign	:	IN STD_LOGIC := '0';
		errdetect	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		fifordin	:	IN STD_LOGIC := '0';
		fifordout	:	OUT STD_LOGIC;
		fiforesetrd	:	IN STD_LOGIC := '0';
		grayelecidleinferselfromtx	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		hip8b10binvpolarity	:	IN STD_LOGIC := '0';
		hipdataout	:	OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		hipdatavalid	:	OUT STD_LOGIC;
		hipelecidle	:	OUT STD_LOGIC;
		hipelecidleinfersel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		hipphydonestatus	:	OUT STD_LOGIC;
		hippowerdown	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		hipstatus	:	OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		invpol	:	IN STD_LOGIC := '0';
		k1detect	:	OUT STD_LOGIC;
		k2detect	:	OUT STD_LOGIC;
		localrefclk	:	IN STD_LOGIC := '0';
		masterclk	:	IN STD_LOGIC := '0';
		parallelfdbk	:	IN STD_LOGIC_VECTOR(19 DOWNTO 0) := (OTHERS => '0');
		patterndetect	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		phfifooverflow	:	OUT STD_LOGIC;
		phfifordenable	:	IN STD_LOGIC := '1';
		phfifordenableout	:	OUT STD_LOGIC;
		phfiforeset	:	IN STD_LOGIC := '0';
		phfiforesetout	:	OUT STD_LOGIC;
		phfifounderflow	:	OUT STD_LOGIC;
		phfifowrdisable	:	IN STD_LOGIC := '0';
		phfifowrdisableout	:	OUT STD_LOGIC;
		phfifox4bytesel	:	IN STD_LOGIC := '0';
		phfifox4rdenable	:	IN STD_LOGIC := '0';
		phfifox4wrclk	:	IN STD_LOGIC := '0';
		phfifox4wrenable	:	IN STD_LOGIC := '0';
		pipe8b10binvpolarity	:	IN STD_LOGIC := '0';
		pipebufferstat	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		pipedatavalid	:	OUT STD_LOGIC;
		pipeelecidle	:	OUT STD_LOGIC;
		pipeenrevparallellpbkfromtx	:	IN STD_LOGIC := '0';
		pipephydonestatus	:	OUT STD_LOGIC;
		pipepowerdown	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		pipepowerstate	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		pipestatetransdoneout	:	OUT STD_LOGIC;
		pipestatus	:	OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		pmatestbusin	:	IN STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		powerdn	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		prbscidenable	:	IN STD_LOGIC := '0';
		quadreset	:	IN STD_LOGIC := '0';
		rdalign	:	OUT STD_LOGIC;
		recoveredclk	:	IN STD_LOGIC := '0';
		refclk	:	IN STD_LOGIC := '0';
		revbitorderwa	:	IN STD_LOGIC := '0';
		revbyteorderwa	:	IN STD_LOGIC := '0';
		revparallelfdbkdata	:	OUT STD_LOGIC_VECTOR(19 DOWNTO 0);
		rlv	:	OUT STD_LOGIC;
		rmfifodatadeleted	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		rmfifodatainserted	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		rmfifoempty	:	OUT STD_LOGIC;
		rmfifofull	:	OUT STD_LOGIC;
		rmfifordena	:	IN STD_LOGIC := '1';
		rmfiforeset	:	IN STD_LOGIC := '0';
		rmfifowrena	:	IN STD_LOGIC := '1';
		runningdisp	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		rxdetectvalid	:	IN STD_LOGIC := '0';
		rxfound	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		signaldetect	:	OUT STD_LOGIC;
		signaldetected	:	IN STD_LOGIC := '0';
		syncstatus	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		syncstatusdeskew	:	OUT STD_LOGIC;
		wareset	:	IN STD_LOGIC := '0';
		xauidelcondmet	:	IN STD_LOGIC := '0';
		xauidelcondmetout	:	OUT STD_LOGIC;
		xauififoovr	:	IN STD_LOGIC := '0';
		xauififoovrout	:	OUT STD_LOGIC;
		xauiinsertincomplete	:	IN STD_LOGIC := '0';
		xauiinsertincompleteout	:	OUT STD_LOGIC;
		xauilatencycomp	:	IN STD_LOGIC := '0';
		xauilatencycompout	:	OUT STD_LOGIC;
		xgmctrldet	:	OUT STD_LOGIC;
		xgmctrlin	:	IN STD_LOGIC := '0';
		xgmdatain	:	IN STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		xgmdataout	:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		xgmdatavalid	:	OUT STD_LOGIC;
		xgmrunningdisp	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneiv_hssi_rx_pma
	 GENERIC 
	 (
		allow_serial_loopback	:	STRING := "false";
		channel_number	:	NATURAL := 0;
		common_mode	:	STRING := "0.82V";
		deserialization_factor	:	NATURAL := 8;
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		effective_data_rate	:	STRING := "UNUSED";
		enable_dpa_shift	:	STRING := "false";
		enable_initial_phase_selection	:	STRING := "true";
		enable_local_divider	:	STRING := "false";
		enable_ltd	:	STRING := "false";
		enable_ltr	:	STRING := "false";
		enable_pd_counter_accumulate_mode	:	STRING := "true";
		enable_second_order_loop	:	STRING := "false";
		eq_dc_gain	:	NATURAL := 0;
		eq_setting	:	NATURAL := 1;
		force_signal_detect	:	STRING := "false";
		initial_phase_value	:	NATURAL := 0;
		logical_channel_address	:	NATURAL := 0;
		loop_1_digital_filter	:	NATURAL := 8;
		offset_cancellation	:	NATURAL := 0;
		pd1_counter_setting	:	NATURAL := 3;
		pd2_counter_setting	:	NATURAL := 2;
		pd_rising_edge_only	:	STRING := "false";
		phase_step_add_setting	:	NATURAL := 2;
		phase_step_sub_setting	:	NATURAL := 1;
		pi_frequency_selector	:	NATURAL := 0;
		ppm_gen1_2_xcnt_en	:	NATURAL := 0;
		ppm_post_eidle	:	NATURAL := 0;
		ppmselect	:	NATURAL := 0;
		protocol_hint	:	STRING := "basic";
		send_reverse_serial_loopback_data	:	STRING := "false";
		send_reverse_serial_loopback_recovered_clk	:	STRING := "false";
		signal_detect_hysteresis	:	NATURAL := 4;
		signal_detect_hysteresis_valid_threshold	:	NATURAL := 14;
		signal_detect_loss_threshold	:	NATURAL := 3;
		termination	:	STRING := "OCT 100 Ohms";
		use_external_termination	:	STRING := "false";
		lpm_type	:	STRING := "cycloneiv_hssi_rx_pma"
	 );
	 PORT
	 ( 
		analogtestbus	:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		clockout	:	OUT STD_LOGIC;
		crupowerdn	:	IN STD_LOGIC := '0';
		datain	:	IN STD_LOGIC := '0';
		datastrobeout	:	OUT STD_LOGIC;
		deserclock	:	IN STD_LOGIC := '0';
		diagnosticlpbkout	:	OUT STD_LOGIC;
		dpashift	:	IN STD_LOGIC := '0';
		dpriodisable	:	IN STD_LOGIC := '1';
		dprioin	:	IN STD_LOGIC_VECTOR(299 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(299 DOWNTO 0);
		freqlocked	:	OUT STD_LOGIC;
		locktodata	:	IN STD_LOGIC := '0';
		locktoref	:	IN STD_LOGIC := '0';
		locktorefout	:	OUT STD_LOGIC;
		powerdn	:	IN STD_LOGIC := '0';
		ppmdetectrefclk	:	IN STD_LOGIC := '0';
		recoverdataout	:	OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		reverselpbkout	:	OUT STD_LOGIC;
		rxpmareset	:	IN STD_LOGIC := '0';
		seriallpbkin	:	IN STD_LOGIC := '0';
		signaldetect	:	OUT STD_LOGIC;
		testbussel	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneiv_hssi_tx_pcs
	 GENERIC 
	 (
		allow_polarity_inversion	:	STRING := "false";
		bitslip_enable	:	STRING := "false";
		channel_bonding	:	STRING := "none";
		channel_number	:	NATURAL := 0;
		channel_width	:	NATURAL := 8;
		core_clock_0ppm	:	STRING := "false";
		datapath_low_latency_mode	:	STRING := "false";
		datapath_protocol	:	STRING := "basic";
		disable_ph_low_latency_mode	:	STRING := "false";
		disparity_mode	:	STRING := "none";
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		elec_idle_delay	:	NATURAL := 3;
		enable_bit_reversal	:	STRING := "false";
		enable_idle_selection	:	STRING := "false";
		enable_phfifo_bypass	:	STRING := "false";
		enable_reverse_parallel_loopback	:	STRING := "false";
		enable_self_test_mode	:	STRING := "false";
		enc_8b_10b_compatibility_mode	:	STRING := "false";
		enc_8b_10b_mode	:	STRING := "none";
		force_echar	:	STRING := "false";
		force_kchar	:	STRING := "false";
		hip_enable	:	STRING := "false";
		logical_channel_address	:	NATURAL := 0;
		ph_fifo_reg_mode	:	STRING := "false";
		ph_fifo_reset_enable	:	STRING := "false";
		ph_fifo_user_ctrl_enable	:	STRING := "false";
		pipe_voltage_swing_control	:	STRING := "false";
		prbs_cid_pattern	:	STRING := "false";
		prbs_cid_pattern_length	:	NATURAL := 0;
		protocol_hint	:	STRING := "basic";
		refclk_select	:	STRING := "local";
		reset_clock_output_during_digital_reset	:	STRING := "false";
		self_test_mode	:	STRING := "crpat";
		use_double_data_mode	:	STRING := "false";
		wr_clk_mux_select	:	STRING := "int_clk";
		lpm_type	:	STRING := "cycloneiv_hssi_tx_pcs"
	 );
	 PORT
	 ( 
		bitslipboundaryselect	:	IN STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
		clkout	:	OUT STD_LOGIC;
		coreclk	:	IN STD_LOGIC := '0';
		coreclkout	:	OUT STD_LOGIC;
		ctrlenable	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		datain	:	IN STD_LOGIC_VECTOR(19 DOWNTO 0) := (OTHERS => '0');
		datainfull	:	IN STD_LOGIC_VECTOR(21 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
		detectrxloop	:	IN STD_LOGIC := '0';
		digitalreset	:	IN STD_LOGIC := '0';
		dispval	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		dpriodisable	:	IN STD_LOGIC := '1';
		dprioin	:	IN STD_LOGIC_VECTOR(149 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(149 DOWNTO 0);
		elecidleinfersel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		enrevparallellpbk	:	IN STD_LOGIC := '0';
		forcedisp	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		forceelecidle	:	IN STD_LOGIC := '0';
		forceelecidleout	:	OUT STD_LOGIC;
		grayelecidleinferselout	:	OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		hipdatain	:	IN STD_LOGIC_VECTOR(9 DOWNTO 0) := (OTHERS => '0');
		hipdetectrxloop	:	IN STD_LOGIC := '0';
		hipelecidleinfersel	:	IN STD_LOGIC_VECTOR(2 DOWNTO 0) := (OTHERS => '0');
		hipforceelecidle	:	IN STD_LOGIC := '0';
		hippowerdn	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		hiptxclkout	:	OUT STD_LOGIC;
		invpol	:	IN STD_LOGIC := '0';
		localrefclk	:	IN STD_LOGIC := '0';
		parallelfdbkout	:	OUT STD_LOGIC_VECTOR(19 DOWNTO 0);
		phfifooverflow	:	OUT STD_LOGIC;
		phfiforddisable	:	IN STD_LOGIC := '0';
		phfiforddisableout	:	OUT STD_LOGIC;
		phfiforeset	:	IN STD_LOGIC := '0';
		phfiforesetout	:	OUT STD_LOGIC;
		phfifounderflow	:	OUT STD_LOGIC;
		phfifowrenable	:	IN STD_LOGIC := '1';
		phfifowrenableout	:	OUT STD_LOGIC;
		phfifox4bytesel	:	IN STD_LOGIC := '0';
		phfifox4rdclk	:	IN STD_LOGIC := '0';
		phfifox4rdenable	:	IN STD_LOGIC := '0';
		phfifox4wrenable	:	IN STD_LOGIC := '0';
		pipeenrevparallellpbkout	:	OUT STD_LOGIC;
		pipepowerdownout	:	OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		pipepowerstateout	:	OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		pipestatetransdone	:	IN STD_LOGIC := '0';
		pipetxswing	:	IN STD_LOGIC := '0';
		powerdn	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0');
		prbscidenable	:	IN STD_LOGIC := '0';
		quadreset	:	IN STD_LOGIC := '0';
		rdenablesync	:	OUT STD_LOGIC;
		refclk	:	IN STD_LOGIC := '0';
		revparallelfdbk	:	IN STD_LOGIC_VECTOR(19 DOWNTO 0) := (OTHERS => '0');
		txdetectrx	:	OUT STD_LOGIC;
		xgmctrl	:	IN STD_LOGIC := '0';
		xgmctrlenable	:	OUT STD_LOGIC;
		xgmdatain	:	IN STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		xgmdataout	:	OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  cycloneiv_hssi_tx_pma
	 GENERIC 
	 (
		channel_number	:	NATURAL := 0;
		common_mode	:	STRING := "0.65V";
		dprio_config_mode	:	STD_LOGIC_VECTOR(5 DOWNTO 0) := "000000";
		effective_data_rate	:	STRING := "UNUSED";
		enable_diagnostic_loopback	:	STRING := "false";
		enable_reverse_serial_loopback	:	STRING := "false";
		enable_txclkout_loopback	:	STRING := "false";
		logical_channel_address	:	NATURAL := 0;
		preemp_tap_1	:	NATURAL := 0;
		protocol_hint	:	STRING := "basic";
		rx_detect	:	NATURAL := 0;
		serialization_factor	:	NATURAL := 8;
		slew_rate	:	STRING := "low";
		termination	:	STRING := "OCT 100 Ohms";
		use_external_termination	:	STRING := "false";
		use_rx_detect	:	STRING := "false";
		vod_selection	:	NATURAL := 0;
		lpm_type	:	STRING := "cycloneiv_hssi_tx_pma"
	 );
	 PORT
	 ( 
		cgbpowerdn	:	IN STD_LOGIC := '0';
		clockout	:	OUT STD_LOGIC;
		datain	:	IN STD_LOGIC_VECTOR(9 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT STD_LOGIC;
		detectrxpowerdown	:	IN STD_LOGIC := '0';
		diagnosticlpbkin	:	IN STD_LOGIC := '0';
		dpriodisable	:	IN STD_LOGIC := '0';
		dprioin	:	IN STD_LOGIC_VECTOR(299 DOWNTO 0) := (OTHERS => '0');
		dprioout	:	OUT STD_LOGIC_VECTOR(299 DOWNTO 0);
		fastrefclk0in	:	IN STD_LOGIC := '0';
		forceelecidle	:	IN STD_LOGIC := '0';
		powerdn	:	IN STD_LOGIC := '0';
		refclk0in	:	IN STD_LOGIC := '0';
		refclk0inpulse	:	IN STD_LOGIC := '0';
		reverselpbkin	:	IN STD_LOGIC := '0';
		rxdetectclk	:	IN STD_LOGIC := '0';
		rxdetecten	:	IN STD_LOGIC := '0';
		rxdetectvalidout	:	OUT STD_LOGIC;
		rxfoundout	:	OUT STD_LOGIC;
		seriallpbkout	:	OUT STD_LOGIC;
		txpmareset	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	wire_w_lg_w_lg_w_lg_fixedclk_sel57w58w59w(0) <= wire_w_lg_w_lg_fixedclk_sel57w58w(0) AND fixedclk_div_in(0);
	wire_w_lg_w_lg_w_lg_fixedclk_sel57w64w65w(0) <= wire_w_lg_w_lg_fixedclk_sel57w64w(0) AND fixedclk_div_in(0);
	wire_w_lg_w_lg_w_lg_fixedclk_sel57w69w70w(0) <= wire_w_lg_w_lg_fixedclk_sel57w69w(0) AND fixedclk_div_in(0);
	wire_w_lg_w_lg_w_lg_fixedclk_sel57w74w75w(0) <= wire_w_lg_w_lg_fixedclk_sel57w74w(0) AND fixedclk_div_in(0);
	wire_w_lg_w_lg_w_lg_fixedclk_sel53w54w55w(0) <= wire_w_lg_w_lg_fixedclk_sel53w54w(0) AND fixedclk;
	wire_w_lg_w_lg_fixedclk_sel57w58w(0) <= wire_w_lg_fixedclk_sel57w(0) AND wire_w_fixedclk_fast_range56w(0);
	wire_w_lg_w_lg_fixedclk_sel57w64w(0) <= wire_w_lg_fixedclk_sel57w(0) AND wire_w_fixedclk_fast_range63w(0);
	wire_w_lg_w_lg_fixedclk_sel57w69w(0) <= wire_w_lg_fixedclk_sel57w(0) AND wire_w_fixedclk_fast_range68w(0);
	wire_w_lg_w_lg_fixedclk_sel57w74w(0) <= wire_w_lg_fixedclk_sel57w(0) AND wire_w_fixedclk_fast_range73w(0);
	wire_w_lg_w_lg_fixedclk_sel53w54w(0) <= wire_w_lg_fixedclk_sel53w(0) AND wire_w_lg_fixedclk_enable52w(0);
	wire_w_lg_w_lg_reconfig_togxb_busy514w515w(0) <= wire_w_lg_reconfig_togxb_busy514w(0) AND wire_w_rx_analogreset_range513w(0);
	wire_w_lg_fixedclk_sel57w(0) <= fixedclk_sel(0) AND fixedclk_enable(0);
	wire_w_lg_fixedclk_enable52w(0) <= NOT fixedclk_enable(0);
	wire_w_lg_fixedclk_sel53w(0) <= NOT fixedclk_sel(0);
	wire_w_lg_reconfig_togxb_busy514w(0) <= NOT reconfig_togxb_busy(0);
	wire_w_lg_w_rx_analogreset_range513w612w(0) <= NOT wire_w_rx_analogreset_range513w(0);
	wire_w_lg_w_lg_w_lg_w_lg_fixedclk_sel57w58w59w60w(0) <= wire_w_lg_w_lg_w_lg_fixedclk_sel57w58w59w(0) OR wire_w_lg_w_lg_w_lg_fixedclk_sel53w54w55w(0);
	wire_w_lg_w_lg_w_lg_w_lg_fixedclk_sel57w64w65w66w(0) <= wire_w_lg_w_lg_w_lg_fixedclk_sel57w64w65w(0) OR wire_w_lg_w_lg_w_lg_fixedclk_sel53w54w55w(0);
	wire_w_lg_w_lg_w_lg_w_lg_fixedclk_sel57w69w70w71w(0) <= wire_w_lg_w_lg_w_lg_fixedclk_sel57w69w70w(0) OR wire_w_lg_w_lg_w_lg_fixedclk_sel53w54w55w(0);
	wire_w_lg_w_lg_w_lg_w_lg_fixedclk_sel57w74w75w76w(0) <= wire_w_lg_w_lg_w_lg_fixedclk_sel57w74w75w(0) OR wire_w_lg_w_lg_w_lg_fixedclk_sel53w54w55w(0);
	cal_blk_powerdown <= '0';
	cent_unit_quadresetout <= ( "000" & wire_cent_unit0_quadresetout);
	cent_unit_rxcrupowerdn <= ( wire_cent_unit0_rxcrupowerdown(3 DOWNTO 0));
	cent_unit_rxibpowerdn <= ( wire_cent_unit0_rxibpowerdown(3 DOWNTO 0));
	cent_unit_rxpcsdprioin <= ( rx_pcsdprioout(1599 DOWNTO 0));
	cent_unit_rxpcsdprioout <= ( wire_cent_unit0_rxpcsdprioout(1599 DOWNTO 0));
	cent_unit_rxpmadprioin <= ( rx_pmadprioout(1199 DOWNTO 0));
	cent_unit_rxpmadprioout <= ( wire_cent_unit0_rxpmadprioout(1199 DOWNTO 0));
	cent_unit_tx_dprioin <= ( tx_txdprioout(599 DOWNTO 0));
	cent_unit_txdetectrxpowerdn <= ( wire_cent_unit0_txdetectrxpowerdown(3 DOWNTO 0));
	cent_unit_txdividerpowerdown <= ( wire_cent_unit0_txdividerpowerdown(3 DOWNTO 0));
	cent_unit_txdprioout <= ( wire_cent_unit0_txpcsdprioout(599 DOWNTO 0));
	cent_unit_txobpowerdn <= ( wire_cent_unit0_txobpowerdown(3 DOWNTO 0));
	cent_unit_txpmadprioin <= ( tx_pmadprioout(1199 DOWNTO 0));
	cent_unit_txpmadprioout <= ( wire_cent_unit0_txpmadprioout(1199 DOWNTO 0));
	coreclkout(0) <= ( coreclkout_wire(0));
	coreclkout_wire(0) <= ( wire_cent_unit0_coreclkout);
	fixedclk_div_in <= fixedclk_div;
	fixedclk_enable(0) <= reconfig_togxb_busy_reg(0);
	fixedclk_fast <= (OTHERS => '1');
	fixedclk_sel(0) <= reconfig_togxb_busy_reg(1);
	fixedclk_to_cmu <= ( wire_w_lg_w_lg_w_lg_w_lg_fixedclk_sel57w74w75w76w & wire_w_lg_w_lg_w_lg_w_lg_fixedclk_sel57w69w70w71w & wire_w_lg_w_lg_w_lg_w_lg_fixedclk_sel57w64w65w66w & wire_w_lg_w_lg_w_lg_w_lg_fixedclk_sel57w58w59w60w);
	hip_tx_clkout <= ( "000" & wire_cent_unit0_refclkout);
	int_pipeenrevparallellpbkfromtx <= ( wire_transmit_pcs3_pipeenrevparallellpbkout & wire_transmit_pcs2_pipeenrevparallellpbkout & wire_transmit_pcs1_pipeenrevparallellpbkout & wire_transmit_pcs0_pipeenrevparallellpbkout);
	int_rx_coreclkout <= ( wire_receive_pcs3_coreclkout & wire_receive_pcs2_coreclkout & wire_receive_pcs1_coreclkout & wire_receive_pcs0_coreclkout);
	int_rx_phfifordenableout <= ( wire_receive_pcs3_phfifordenableout & wire_receive_pcs2_phfifordenableout & wire_receive_pcs1_phfifordenableout & wire_receive_pcs0_phfifordenableout);
	int_rx_phfiforesetout <= ( wire_receive_pcs3_phfiforesetout & wire_receive_pcs2_phfiforesetout & wire_receive_pcs1_phfiforesetout & wire_receive_pcs0_phfiforesetout);
	int_rx_phfifowrdisableout <= ( wire_receive_pcs3_phfifowrdisableout & wire_receive_pcs2_phfifowrdisableout & wire_receive_pcs1_phfifowrdisableout & wire_receive_pcs0_phfifowrdisableout);
	int_rx_phfifoxnbytesel <= ( int_rxphfifox4byteselout(0) & int_rxphfifox4byteselout(0) & int_rxphfifox4byteselout(0) & int_rxphfifox4byteselout(0));
	int_rx_phfifoxnrdenable <= ( int_rxphfifox4rdenableout(0) & int_rxphfifox4rdenableout(0) & int_rxphfifox4rdenableout(0) & int_rxphfifox4rdenableout(0));
	int_rx_phfifoxnwrclk <= ( int_rxphfifox4wrclkout(0) & int_rxphfifox4wrclkout(0) & int_rxphfifox4wrclkout(0) & int_rxphfifox4wrclkout(0));
	int_rx_phfifoxnwrenable <= ( int_rxphfifox4wrenableout(0) & int_rxphfifox4wrenableout(0) & int_rxphfifox4wrenableout(0) & int_rxphfifox4wrenableout(0));
	int_rxcoreclk(0) <= ( int_rx_coreclkout(0));
	int_rxphfifordenable(0) <= ( int_rx_phfifordenableout(0));
	int_rxphfiforeset(0) <= ( int_rx_phfiforesetout(0));
	int_rxphfifox4byteselout(0) <= ( wire_cent_unit0_rxphfifox4byteselout);
	int_rxphfifox4rdenableout(0) <= ( wire_cent_unit0_rxphfifox4rdenableout);
	int_rxphfifox4wrclkout(0) <= ( wire_cent_unit0_rxphfifox4wrclkout);
	int_rxphfifox4wrenableout(0) <= ( wire_cent_unit0_rxphfifox4wrenableout);
	int_tx_coreclkout <= ( wire_transmit_pcs3_coreclkout & wire_transmit_pcs2_coreclkout & wire_transmit_pcs1_coreclkout & wire_transmit_pcs0_coreclkout);
	int_tx_phfiforddisableout <= ( wire_transmit_pcs3_phfiforddisableout & wire_transmit_pcs2_phfiforddisableout & wire_transmit_pcs1_phfiforddisableout & wire_transmit_pcs0_phfiforddisableout);
	int_tx_phfiforesetout <= ( wire_transmit_pcs3_phfiforesetout & wire_transmit_pcs2_phfiforesetout & wire_transmit_pcs1_phfiforesetout & wire_transmit_pcs0_phfiforesetout);
	int_tx_phfifowrenableout <= ( wire_transmit_pcs3_phfifowrenableout & wire_transmit_pcs2_phfifowrenableout & wire_transmit_pcs1_phfifowrenableout & wire_transmit_pcs0_phfifowrenableout);
	int_tx_phfifoxnbytesel <= ( int_txphfifox4byteselout(0) & int_txphfifox4byteselout(0) & int_txphfifox4byteselout(0) & int_txphfifox4byteselout(0));
	int_tx_phfifoxnrdclk <= ( int_txphfifox4rdclkout(0) & int_txphfifox4rdclkout(0) & int_txphfifox4rdclkout(0) & int_txphfifox4rdclkout(0));
	int_tx_phfifoxnrdenable <= ( int_txphfifox4rdenableout(0) & int_txphfifox4rdenableout(0) & int_txphfifox4rdenableout(0) & int_txphfifox4rdenableout(0));
	int_tx_phfifoxnwrenable <= ( int_txphfifox4wrenableout(0) & int_txphfifox4wrenableout(0) & int_txphfifox4wrenableout(0) & int_txphfifox4wrenableout(0));
	int_txcoreclk(0) <= ( int_tx_coreclkout(0));
	int_txphfiforddisable(0) <= ( int_tx_phfiforddisableout(0));
	int_txphfiforeset(0) <= ( int_tx_phfiforesetout(0));
	int_txphfifowrenable(0) <= ( int_tx_phfifowrenableout(0));
	int_txphfifox4byteselout(0) <= ( wire_cent_unit0_txphfifox4byteselout);
	int_txphfifox4rdclkout(0) <= ( wire_cent_unit0_txphfifox4rdclkout);
	int_txphfifox4rdenableout(0) <= ( wire_cent_unit0_txphfifox4rdenableout);
	int_txphfifox4wrenableout(0) <= ( wire_cent_unit0_txphfifox4wrenableout);
	nonusertocmu_out(0) <= ( wire_cal_blk0_nonusertocmu);
	pipedatavalid <= ( pipedatavalid_out(3 DOWNTO 0));
	pipedatavalid_out <= ( wire_receive_pcs3_hipdatavalid & wire_receive_pcs2_hipdatavalid & wire_receive_pcs1_hipdatavalid & wire_receive_pcs0_hipdatavalid);
	pipeelecidle <= ( pipeelecidle_out(3 DOWNTO 0));
	pipeelecidle_out <= ( wire_receive_pcs3_hipelecidle & wire_receive_pcs2_hipelecidle & wire_receive_pcs1_hipelecidle & wire_receive_pcs0_hipelecidle);
	pipephydonestatus <= ( wire_receive_pcs3_hipphydonestatus & wire_receive_pcs2_hipphydonestatus & wire_receive_pcs1_hipphydonestatus & wire_receive_pcs0_hipphydonestatus);
	pipestatus <= ( wire_receive_pcs3_hipstatus & wire_receive_pcs2_hipstatus & wire_receive_pcs1_hipstatus & wire_receive_pcs0_hipstatus);
	pll_locked(0) <= ( wire_pll0_locked);
	pll_powerdown <= (OTHERS => '0');
	reconfig_fromgxb <= ( rx_pma_analogtestbus(4 DOWNTO 1) & wire_cent_unit0_dprioout);
	reconfig_togxb_busy(0) <= reconfig_togxb(3);
	reconfig_togxb_disable(0) <= reconfig_togxb(1);
	reconfig_togxb_in(0) <= reconfig_togxb(0);
	reconfig_togxb_load(0) <= reconfig_togxb(2);
	refclk_pma(0) <= ( wire_cent_unit0_refclkout);
	rx_analogreset_in <= ( wire_w_lg_w_lg_reconfig_togxb_busy514w515w & wire_w_lg_w_lg_reconfig_togxb_busy514w515w & wire_w_lg_w_lg_reconfig_togxb_busy514w515w & wire_w_lg_w_lg_reconfig_togxb_busy514w515w);
	rx_analogreset_out <= ( wire_cent_unit0_rxanalogresetout(3 DOWNTO 0));
	rx_ctrldetect <= ( wire_receive_pcs3_hipdataout(8) & wire_receive_pcs2_hipdataout(8) & wire_receive_pcs1_hipdataout(8) & wire_receive_pcs0_hipdataout(8));
	rx_dataout <= ( rx_out_wire(31 DOWNTO 0));
	rx_deserclock_in <= ( wire_pll0_icdrclk & wire_pll0_icdrclk & wire_pll0_icdrclk & wire_pll0_icdrclk);
	rx_digitalreset_in <= ( rx_digitalreset(0) & rx_digitalreset(0) & rx_digitalreset(0) & rx_digitalreset(0));
	rx_digitalreset_out <= ( wire_cent_unit0_rxdigitalresetout(3 DOWNTO 0));
	rx_enapatternalign <= (OTHERS => '0');
	rx_freqlocked <= ( wire_receive_pma3_w_lg_freqlocked815w & wire_receive_pma2_w_lg_freqlocked748w & wire_receive_pma1_w_lg_freqlocked681w & wire_receive_pma0_w_lg_freqlocked613w);
	rx_locktodata <= (OTHERS => '0');
	rx_locktorefclk_wire <= ( wire_receive_pcs3_cdrctrllocktorefclkout & wire_receive_pcs2_cdrctrllocktorefclkout & wire_receive_pcs1_cdrctrllocktorefclkout & wire_receive_pcs0_cdrctrllocktorefclkout);
	rx_out_wire <= ( wire_receive_pcs3_hipdataout(7 DOWNTO 0) & wire_receive_pcs2_hipdataout(7 DOWNTO 0) & wire_receive_pcs1_hipdataout(7 DOWNTO 0) & wire_receive_pcs0_hipdataout(7 DOWNTO 0));
	rx_pcs_rxfound_wire <= ( txdetectrxout(3) & tx_rxfoundout(3) & txdetectrxout(2) & tx_rxfoundout(2) & txdetectrxout(1) & tx_rxfoundout(1) & txdetectrxout(0) & tx_rxfoundout(0));
	rx_pcsdprioin_wire <= ( cent_unit_rxpcsdprioout(1599 DOWNTO 0));
	rx_pcsdprioout <= ( wire_receive_pcs3_dprioout & wire_receive_pcs2_dprioout & wire_receive_pcs1_dprioout & wire_receive_pcs0_dprioout);
	rx_phfifordenable <= (OTHERS => '1');
	rx_phfiforeset <= (OTHERS => '0');
	rx_phfifowrdisable <= (OTHERS => '0');
	rx_pll_pfdrefclkout_wire <= ( wire_pll0_fref & wire_pll0_fref & wire_pll0_fref & wire_pll0_fref);
	rx_pma_analogtestbus <= ( "0" & wire_receive_pma3_analogtestbus(6) & wire_receive_pma2_analogtestbus(6) & wire_receive_pma1_analogtestbus(6) & wire_receive_pma0_analogtestbus(6));
	rx_pma_clockout <= ( wire_receive_pma3_clockout & wire_receive_pma2_clockout & wire_receive_pma1_clockout & wire_receive_pma0_clockout);
	rx_pma_recoverdataout_wire <= ( wire_receive_pma3_recoverdataout(9 DOWNTO 0) & wire_receive_pma2_recoverdataout(9 DOWNTO 0) & wire_receive_pma1_recoverdataout(9 DOWNTO 0) & wire_receive_pma0_recoverdataout(9 DOWNTO 0));
	rx_pmadprioin_wire <= ( cent_unit_rxpmadprioout(1199 DOWNTO 0));
	rx_pmadprioout <= ( wire_receive_pma3_dprioout & wire_receive_pma2_dprioout & wire_receive_pma1_dprioout & wire_receive_pma0_dprioout);
	rx_powerdown <= (OTHERS => '0');
	rx_powerdown_in <= ( rx_powerdown(3 DOWNTO 0));
	rx_prbscidenable <= (OTHERS => '0');
	rx_reverselpbkout <= ( wire_receive_pma3_reverselpbkout & wire_receive_pma2_reverselpbkout & wire_receive_pma1_reverselpbkout & wire_receive_pma0_reverselpbkout);
	rx_revparallelfdbkdata <= ( wire_receive_pcs3_revparallelfdbkdata & wire_receive_pcs2_revparallelfdbkdata & wire_receive_pcs1_revparallelfdbkdata & wire_receive_pcs0_revparallelfdbkdata);
	rx_rmfiforeset <= (OTHERS => '0');
	rx_signaldetect_wire <= ( wire_receive_pma3_signaldetect & wire_receive_pma2_signaldetect & wire_receive_pma1_signaldetect & wire_receive_pma0_signaldetect);
	rxphfifowrdisable(0) <= ( int_rx_phfifowrdisableout(0));
	tx_analogreset_out <= ( wire_cent_unit0_txanalogresetout(3 DOWNTO 0));
	tx_datain_wire <= ( tx_datain(31 DOWNTO 0));
	tx_dataout <= ( txdataout(3 DOWNTO 0));
	tx_dataout_pcs_to_pma <= ( wire_transmit_pcs3_dataout(9 DOWNTO 0) & wire_transmit_pcs2_dataout(9 DOWNTO 0) & wire_transmit_pcs1_dataout(9 DOWNTO 0) & wire_transmit_pcs0_dataout(9 DOWNTO 0));
	tx_diagnosticlpbkin <= ( wire_receive_pma3_diagnosticlpbkout & wire_receive_pma2_diagnosticlpbkout & wire_receive_pma1_diagnosticlpbkout & wire_receive_pma0_diagnosticlpbkout);
	tx_digitalreset_in <= ( tx_digitalreset(0) & tx_digitalreset(0) & tx_digitalreset(0) & tx_digitalreset(0));
	tx_digitalreset_out <= ( wire_cent_unit0_txdigitalresetout(3 DOWNTO 0));
	tx_dprioin_wire <= ( cent_unit_txdprioout(599 DOWNTO 0));
	tx_invpolarity <= (OTHERS => '0');
	tx_localrefclk <= ( wire_transmit_pma3_clockout & wire_transmit_pma2_clockout & wire_transmit_pma1_clockout & wire_transmit_pma0_clockout);
	tx_pcs_forceelecidleout <= ( wire_transmit_pcs3_forceelecidleout & wire_transmit_pcs2_forceelecidleout & wire_transmit_pcs1_forceelecidleout & wire_transmit_pcs0_forceelecidleout);
	tx_phfiforeset <= (OTHERS => '0');
	tx_pipepowerdownout <= ( wire_transmit_pcs3_pipepowerdownout & wire_transmit_pcs2_pipepowerdownout & wire_transmit_pcs1_pipepowerdownout & wire_transmit_pcs0_pipepowerdownout);
	tx_pipepowerstateout <= ( wire_transmit_pcs3_pipepowerstateout & wire_transmit_pcs2_pipepowerstateout & wire_transmit_pcs1_pipepowerstateout & wire_transmit_pcs0_pipepowerstateout);
	tx_pma_fastrefclk0in <= ( wire_pll0_clk(0) & wire_pll0_clk(0) & wire_pll0_clk(0) & wire_pll0_clk(0));
	tx_pma_refclk0in <= ( wire_pll0_clk(1) & wire_pll0_clk(1) & wire_pll0_clk(1) & wire_pll0_clk(1));
	tx_pma_refclk0inpulse <= ( wire_pll0_clk(2) & wire_pll0_clk(2) & wire_pll0_clk(2) & wire_pll0_clk(2));
	tx_pmadprioin_wire <= ( cent_unit_txpmadprioout(1199 DOWNTO 0));
	tx_pmadprioout <= ( wire_transmit_pma3_dprioout & wire_transmit_pma2_dprioout & wire_transmit_pma1_dprioout & wire_transmit_pma0_dprioout);
	tx_revparallellpbken <= (OTHERS => '0');
	tx_rxdetectvalidout <= ( wire_transmit_pma3_rxdetectvalidout & wire_transmit_pma2_rxdetectvalidout & wire_transmit_pma1_rxdetectvalidout & wire_transmit_pma0_rxdetectvalidout);
	tx_rxfoundout <= ( wire_transmit_pma3_rxfoundout & wire_transmit_pma2_rxfoundout & wire_transmit_pma1_rxfoundout & wire_transmit_pma0_rxfoundout);
	tx_serialloopbackout <= ( wire_transmit_pma3_seriallpbkout & wire_transmit_pma2_seriallpbkout & wire_transmit_pma1_seriallpbkout & wire_transmit_pma0_seriallpbkout);
	tx_txdprioout <= ( wire_transmit_pcs3_dprioout & wire_transmit_pcs2_dprioout & wire_transmit_pcs1_dprioout & wire_transmit_pcs0_dprioout);
	txdataout <= ( wire_transmit_pma3_dataout & wire_transmit_pma2_dataout & wire_transmit_pma1_dataout & wire_transmit_pma0_dataout);
	txdetectrxout <= ( wire_transmit_pcs3_txdetectrx & wire_transmit_pcs2_txdetectrx & wire_transmit_pcs1_txdetectrx & wire_transmit_pcs0_txdetectrx);
	w_cent_unit_dpriodisableout1w(0) <= ( wire_cent_unit0_dpriodisableout);
	wire_w_fixedclk_fast_range56w(0) <= fixedclk_fast(0);
	wire_w_fixedclk_fast_range63w(0) <= fixedclk_fast(1);
	wire_w_fixedclk_fast_range68w(0) <= fixedclk_fast(2);
	wire_w_fixedclk_fast_range73w(0) <= fixedclk_fast(3);
	wire_w_rx_analogreset_range513w(0) <= rx_analogreset(0);
	wire_pll0_areset <= wire_w_lg_w_pll_areset_range50w51w(0);
	wire_w_lg_w_pll_areset_range50w51w(0) <= pll_areset(0) OR pll_powerdown(0);
	wire_pll0_inclk <= ( "0" & pll_inclk(0));
	pll0 :  altpll
	  GENERIC MAP (
		bandwidth_type => "AUTO",
		clk0_divide_by => 2,
		clk0_multiply_by => 25,
		clk1_divide_by => 10,
		clk1_multiply_by => 25,
		clk2_divide_by => 10,
		clk2_duty_cycle => 20,
		clk2_multiply_by => 25,
		DPA_DIVIDE_BY => 2,
		DPA_MULTIPLY_BY => 25,
		inclk0_input_frequency => 10000,
		operation_mode => "no_compensation",
		INTENDED_DEVICE_FAMILY => "Cyclone IV GX"
	  )
	  PORT MAP ( 
		areset => wire_pll0_areset,
		clk => wire_pll0_clk,
		fref => wire_pll0_fref,
		icdrclk => wire_pll0_icdrclk,
		inclk => wire_pll0_inclk,
		locked => wire_pll0_locked
	  );
	cal_blk0 :  cycloneiv_hssi_calibration_block
	  PORT MAP ( 
		clk => cal_blk_clk,
		nonusertocmu => wire_cal_blk0_nonusertocmu,
		powerdn => cal_blk_powerdown
	  );
	wire_cent_unit0_adet <= (OTHERS => '0');
	wire_cent_unit0_fixedclk <= ( fixedclk_to_cmu(3 DOWNTO 0));
	wire_cent_unit0_rdalign <= (OTHERS => '0');
	wire_cent_unit0_rxanalogreset <= ( rx_analogreset_in(3 DOWNTO 0));
	wire_cent_unit0_rxctrl <= (OTHERS => '0');
	wire_cent_unit0_rxdatain <= (OTHERS => '0');
	wire_cent_unit0_rxdatavalid <= (OTHERS => '0');
	wire_cent_unit0_rxdigitalreset <= ( rx_digitalreset_in(3 DOWNTO 0));
	wire_cent_unit0_rxpcsdprioin <= ( cent_unit_rxpcsdprioin(1599 DOWNTO 0));
	wire_cent_unit0_rxpmadprioin <= ( cent_unit_rxpmadprioin(1199 DOWNTO 0));
	wire_cent_unit0_rxpowerdown <= ( rx_powerdown_in(3 DOWNTO 0));
	wire_cent_unit0_rxrunningdisp <= (OTHERS => '0');
	wire_cent_unit0_syncstatus <= (OTHERS => '0');
	wire_cent_unit0_txctrl <= (OTHERS => '0');
	wire_cent_unit0_txdatain <= (OTHERS => '0');
	wire_cent_unit0_txdigitalreset <= ( tx_digitalreset_in(3 DOWNTO 0));
	wire_cent_unit0_txpcsdprioin <= ( cent_unit_tx_dprioin(599 DOWNTO 0));
	wire_cent_unit0_txpmadprioin <= ( cent_unit_txpmadprioin(1199 DOWNTO 0));
	cent_unit0 :  cycloneiv_hssi_cmu
	  GENERIC MAP (
		auto_spd_deassert_ph_fifo_rst_count => 8,
		auto_spd_phystatus_notify_count => 14,
		devaddr => ((((starting_channel_number / 4) + 0) MOD 32) + 1),
		dprio_config_mode => "000001",
		in_xaui_mode => "false",
		portaddr => (((starting_channel_number + 0) / 128) + 1),
		rx0_channel_bonding => "x4",
		rx0_clk1_mux_select => "recovered clock",
		rx0_clk2_mux_select => "digital reference clock",
		rx0_ph_fifo_reg_mode => "true",
		rx0_rd_clk_mux_select => "int clock",
		rx0_recovered_clk_mux_select => "recovered clock",
		rx0_reset_clock_output_during_digital_reset => "false",
		rx0_use_double_data_mode => "false",
		tx0_channel_bonding => "x4",
		tx0_rd_clk_mux_select => "central",
		tx0_reset_clock_output_during_digital_reset => "false",
		tx0_use_double_data_mode => "false",
		tx0_wr_clk_mux_select => "int_clk",
		use_coreclk_out_post_divider => "false",
		use_deskew_fifo => "false"
	  )
	  PORT MAP ( 
		adet => wire_cent_unit0_adet,
		coreclkout => wire_cent_unit0_coreclkout,
		dpclk => reconfig_clk,
		dpriodisable => reconfig_togxb_disable(0),
		dpriodisableout => wire_cent_unit0_dpriodisableout,
		dprioin => reconfig_togxb_in(0),
		dprioload => reconfig_togxb_load(0),
		dprioout => wire_cent_unit0_dprioout,
		fixedclk => wire_cent_unit0_fixedclk,
		nonuserfromcal => nonusertocmu_out(0),
		quadreset => gxb_powerdown(0),
		quadresetout => wire_cent_unit0_quadresetout,
		rdalign => wire_cent_unit0_rdalign,
		rdenablesync => wire_gnd,
		recovclk => wire_gnd,
		refclkout => wire_cent_unit0_refclkout,
		rxanalogreset => wire_cent_unit0_rxanalogreset,
		rxanalogresetout => wire_cent_unit0_rxanalogresetout,
		rxcoreclk => int_rxcoreclk(0),
		rxcrupowerdown => wire_cent_unit0_rxcrupowerdown,
		rxctrl => wire_cent_unit0_rxctrl,
		rxdatain => wire_cent_unit0_rxdatain,
		rxdatavalid => wire_cent_unit0_rxdatavalid,
		rxdigitalreset => wire_cent_unit0_rxdigitalreset,
		rxdigitalresetout => wire_cent_unit0_rxdigitalresetout,
		rxibpowerdown => wire_cent_unit0_rxibpowerdown,
		rxpcsdprioin => wire_cent_unit0_rxpcsdprioin,
		rxpcsdprioout => wire_cent_unit0_rxpcsdprioout,
		rxphfifordenable => int_rxphfifordenable(0),
		rxphfiforeset => int_rxphfiforeset(0),
		rxphfifowrdisable => rxphfifowrdisable(0),
		rxphfifox4byteselout => wire_cent_unit0_rxphfifox4byteselout,
		rxphfifox4rdenableout => wire_cent_unit0_rxphfifox4rdenableout,
		rxphfifox4wrclkout => wire_cent_unit0_rxphfifox4wrclkout,
		rxphfifox4wrenableout => wire_cent_unit0_rxphfifox4wrenableout,
		rxpmadprioin => wire_cent_unit0_rxpmadprioin,
		rxpmadprioout => wire_cent_unit0_rxpmadprioout,
		rxpowerdown => wire_cent_unit0_rxpowerdown,
		rxrunningdisp => wire_cent_unit0_rxrunningdisp,
		syncstatus => wire_cent_unit0_syncstatus,
		txanalogresetout => wire_cent_unit0_txanalogresetout,
		txclk => tx_localrefclk(0),
		txcoreclk => int_txcoreclk(0),
		txctrl => wire_cent_unit0_txctrl,
		txdatain => wire_cent_unit0_txdatain,
		txdetectrxpowerdown => wire_cent_unit0_txdetectrxpowerdown,
		txdigitalreset => wire_cent_unit0_txdigitalreset,
		txdigitalresetout => wire_cent_unit0_txdigitalresetout,
		txdividerpowerdown => wire_cent_unit0_txdividerpowerdown,
		txobpowerdown => wire_cent_unit0_txobpowerdown,
		txpcsdprioin => wire_cent_unit0_txpcsdprioin,
		txpcsdprioout => wire_cent_unit0_txpcsdprioout,
		txphfiforddisable => int_txphfiforddisable(0),
		txphfiforeset => int_txphfiforeset(0),
		txphfifowrenable => int_txphfifowrenable(0),
		txphfifox4byteselout => wire_cent_unit0_txphfifox4byteselout,
		txphfifox4rdclkout => wire_cent_unit0_txphfifox4rdclkout,
		txphfifox4rdenableout => wire_cent_unit0_txphfifox4rdenableout,
		txphfifox4wrenableout => wire_cent_unit0_txphfifox4wrenableout,
		txpmadprioin => wire_cent_unit0_txpmadprioin,
		txpmadprioout => wire_cent_unit0_txpmadprioout
	  );
	wire_receive_pcs0_hipelecidleinfersel <= (OTHERS => '0');
	wire_receive_pcs0_parallelfdbk <= (OTHERS => '0');
	wire_receive_pcs0_xgmdatain <= (OTHERS => '0');
	receive_pcs0 :  cycloneiv_hssi_rx_pcs
	  GENERIC MAP (
		align_pattern => "0101111100",
		align_pattern_length => 10,
		allow_align_polarity_inversion => "false",
		allow_pipe_polarity_inversion => "true",
		auto_spd_deassert_ph_fifo_rst_count => 8,
		auto_spd_phystatus_notify_count => 14,
		bit_slip_enable => "false",
		byte_order_invalid_code_or_run_disp_error => "true",
		byte_order_mode => "none",
		byte_order_pad_pattern => "0",
		byte_order_pattern => "0",
		byte_order_pld_ctrl_enable => "false",
		cdrctrl_bypass_ppm_detector_cycle => 1000,
		cdrctrl_cid_mode_enable => "true",
		cdrctrl_enable => "true",
		cdrctrl_mask_cycle => 800,
		cdrctrl_min_lock_to_ref_cycle => 63,
		cdrctrl_rxvalid_mask => "true",
		channel_bonding => "x4",
		channel_number => ((starting_channel_number + 0) MOD 4),
		channel_width => 8,
		clk1_mux_select => "recovered clock",
		clk2_mux_select => "digital reference clock",
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "pipe",
		dec_8b_10b_compatibility_mode => "true",
		dec_8b_10b_mode => "normal",
		deskew_pattern => "0",
		disable_auto_idle_insertion => "false",
		disable_running_disp_in_word_align => "false",
		disallow_kchar_after_pattern_ordered_set => "false",
		dprio_config_mode => "000001",
		elec_idle_gen1_sigdet_enable => "true",
		elec_idle_infer_enable => "false",
		elec_idle_num_com_detect => 3,
		enable_bit_reversal => "false",
		enable_self_test_mode => "false",
		force_signal_detect_dig => "true",
		hip_enable => "true",
		infiniband_invalid_code => 0,
		insert_pad_on_underflow => "false",
		num_align_code_groups_in_ordered_set => 0,
		num_align_cons_good_data => 16,
		num_align_cons_pat => 4,
		num_align_loss_sync_error => 17,
		ph_fifo_low_latency_enable => "true",
		ph_fifo_reg_mode => "true",
		protocol_hint => "pcie",
		rate_match_back_to_back => "false",
		rate_match_delete_threshold => 13,
		rate_match_empty_threshold => 5,
		rate_match_fifo_mode => "true",
		rate_match_full_threshold => 20,
		rate_match_insert_threshold => 11,
		rate_match_ordered_set_based => "false",
		rate_match_pattern1 => "11010000111010000011",
		rate_match_pattern2 => "00101111000101111100",
		rate_match_pattern_size => 20,
		rate_match_pipe_enable => "true",
		rate_match_reset_enable => "false",
		rate_match_skip_set_based => "true",
		rate_match_start_threshold => 7,
		rd_clk_mux_select => "int clock",
		recovered_clk_mux_select => "recovered clock",
		run_length => 40,
		run_length_enable => "true",
		rx_detect_bypass => "false",
		rx_phfifo_wait_cnt => 32,
		rxstatus_error_report_mode => 1,
		self_test_mode => "incremental",
		use_alignment_state_machine => "true",
		use_deskew_fifo => "false",
		use_double_data_mode => "false",
		use_parallel_loopback => "false"
	  )
	  PORT MAP ( 
		a1a2size => wire_gnd,
		alignstatus => wire_gnd,
		alignstatussync => wire_gnd,
		cdrctrlearlyeios => wire_receive_pcs0_cdrctrlearlyeios,
		cdrctrllocktorefclkout => wire_receive_pcs0_cdrctrllocktorefclkout,
		coreclkout => wire_receive_pcs0_coreclkout,
		datain => rx_pma_recoverdataout_wire(9 DOWNTO 0),
		digitalreset => rx_digitalreset_out(0),
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => rx_pcsdprioin_wire(399 DOWNTO 0),
		dprioout => wire_receive_pcs0_dprioout,
		enabledeskew => wire_gnd,
		enabyteord => wire_gnd,
		enapatternalign => rx_enapatternalign(0),
		fifordin => wire_gnd,
		fiforesetrd => wire_gnd,
		hip8b10binvpolarity => pipe8b10binvpolarity(0),
		hipdataout => wire_receive_pcs0_hipdataout,
		hipdatavalid => wire_receive_pcs0_hipdatavalid,
		hipelecidle => wire_receive_pcs0_hipelecidle,
		hipelecidleinfersel => wire_receive_pcs0_hipelecidleinfersel,
		hipphydonestatus => wire_receive_pcs0_hipphydonestatus,
		hippowerdown => powerdn(1 DOWNTO 0),
		hipstatus => wire_receive_pcs0_hipstatus,
		invpol => wire_gnd,
		localrefclk => tx_localrefclk(0),
		masterclk => wire_gnd,
		parallelfdbk => wire_receive_pcs0_parallelfdbk,
		phfifordenable => rx_phfifordenable(0),
		phfifordenableout => wire_receive_pcs0_phfifordenableout,
		phfiforeset => rx_phfiforeset(0),
		phfiforesetout => wire_receive_pcs0_phfiforesetout,
		phfifowrdisable => rx_phfifowrdisable(0),
		phfifowrdisableout => wire_receive_pcs0_phfifowrdisableout,
		phfifox4bytesel => int_rx_phfifoxnbytesel(0),
		phfifox4rdenable => int_rx_phfifoxnrdenable(0),
		phfifox4wrclk => int_rx_phfifoxnwrclk(0),
		phfifox4wrenable => int_rx_phfifoxnwrenable(0),
		pipeenrevparallellpbkfromtx => int_pipeenrevparallellpbkfromtx(0),
		pipepowerdown => tx_pipepowerdownout(1 DOWNTO 0),
		pipepowerstate => tx_pipepowerstateout(3 DOWNTO 0),
		prbscidenable => rx_prbscidenable(0),
		quadreset => cent_unit_quadresetout(0),
		recoveredclk => rx_pma_clockout(0),
		refclk => refclk_pma(0),
		revbitorderwa => wire_gnd,
		revparallelfdbkdata => wire_receive_pcs0_revparallelfdbkdata,
		rmfifordena => wire_gnd,
		rmfiforeset => rx_rmfiforeset(0),
		rmfifowrena => wire_gnd,
		rxdetectvalid => tx_rxdetectvalidout(0),
		rxfound => rx_pcs_rxfound_wire(1 DOWNTO 0),
		signaldetected => rx_signaldetect_wire(0),
		xgmctrlin => wire_gnd,
		xgmdatain => wire_receive_pcs0_xgmdatain
	  );
	wire_receive_pcs1_hipelecidleinfersel <= (OTHERS => '0');
	wire_receive_pcs1_parallelfdbk <= (OTHERS => '0');
	wire_receive_pcs1_xgmdatain <= (OTHERS => '0');
	receive_pcs1 :  cycloneiv_hssi_rx_pcs
	  GENERIC MAP (
		align_pattern => "0101111100",
		align_pattern_length => 10,
		allow_align_polarity_inversion => "false",
		allow_pipe_polarity_inversion => "true",
		auto_spd_deassert_ph_fifo_rst_count => 8,
		auto_spd_phystatus_notify_count => 14,
		bit_slip_enable => "false",
		byte_order_invalid_code_or_run_disp_error => "true",
		byte_order_mode => "none",
		byte_order_pad_pattern => "0",
		byte_order_pattern => "0",
		byte_order_pld_ctrl_enable => "false",
		cdrctrl_bypass_ppm_detector_cycle => 1000,
		cdrctrl_cid_mode_enable => "true",
		cdrctrl_enable => "true",
		cdrctrl_mask_cycle => 800,
		cdrctrl_min_lock_to_ref_cycle => 63,
		cdrctrl_rxvalid_mask => "true",
		channel_bonding => "x4",
		channel_number => ((starting_channel_number + 1) MOD 4),
		channel_width => 8,
		clk1_mux_select => "recovered clock",
		clk2_mux_select => "digital reference clock",
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "pipe",
		dec_8b_10b_compatibility_mode => "true",
		dec_8b_10b_mode => "normal",
		deskew_pattern => "0",
		disable_auto_idle_insertion => "false",
		disable_running_disp_in_word_align => "false",
		disallow_kchar_after_pattern_ordered_set => "false",
		dprio_config_mode => "000001",
		elec_idle_gen1_sigdet_enable => "true",
		elec_idle_infer_enable => "false",
		elec_idle_num_com_detect => 3,
		enable_bit_reversal => "false",
		enable_self_test_mode => "false",
		force_signal_detect_dig => "true",
		hip_enable => "true",
		infiniband_invalid_code => 0,
		insert_pad_on_underflow => "false",
		num_align_code_groups_in_ordered_set => 0,
		num_align_cons_good_data => 16,
		num_align_cons_pat => 4,
		num_align_loss_sync_error => 17,
		ph_fifo_low_latency_enable => "true",
		ph_fifo_reg_mode => "true",
		protocol_hint => "pcie",
		rate_match_back_to_back => "false",
		rate_match_delete_threshold => 13,
		rate_match_empty_threshold => 5,
		rate_match_fifo_mode => "true",
		rate_match_full_threshold => 20,
		rate_match_insert_threshold => 11,
		rate_match_ordered_set_based => "false",
		rate_match_pattern1 => "11010000111010000011",
		rate_match_pattern2 => "00101111000101111100",
		rate_match_pattern_size => 20,
		rate_match_pipe_enable => "true",
		rate_match_reset_enable => "false",
		rate_match_skip_set_based => "true",
		rate_match_start_threshold => 7,
		rd_clk_mux_select => "int clock",
		recovered_clk_mux_select => "recovered clock",
		run_length => 40,
		run_length_enable => "true",
		rx_detect_bypass => "false",
		rx_phfifo_wait_cnt => 32,
		rxstatus_error_report_mode => 1,
		self_test_mode => "incremental",
		use_alignment_state_machine => "true",
		use_deskew_fifo => "false",
		use_double_data_mode => "false",
		use_parallel_loopback => "false"
	  )
	  PORT MAP ( 
		a1a2size => wire_gnd,
		alignstatus => wire_gnd,
		alignstatussync => wire_gnd,
		cdrctrlearlyeios => wire_receive_pcs1_cdrctrlearlyeios,
		cdrctrllocktorefclkout => wire_receive_pcs1_cdrctrllocktorefclkout,
		coreclkout => wire_receive_pcs1_coreclkout,
		datain => rx_pma_recoverdataout_wire(19 DOWNTO 10),
		digitalreset => rx_digitalreset_out(1),
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => rx_pcsdprioin_wire(799 DOWNTO 400),
		dprioout => wire_receive_pcs1_dprioout,
		enabledeskew => wire_gnd,
		enabyteord => wire_gnd,
		enapatternalign => rx_enapatternalign(1),
		fifordin => wire_gnd,
		fiforesetrd => wire_gnd,
		hip8b10binvpolarity => pipe8b10binvpolarity(1),
		hipdataout => wire_receive_pcs1_hipdataout,
		hipdatavalid => wire_receive_pcs1_hipdatavalid,
		hipelecidle => wire_receive_pcs1_hipelecidle,
		hipelecidleinfersel => wire_receive_pcs1_hipelecidleinfersel,
		hipphydonestatus => wire_receive_pcs1_hipphydonestatus,
		hippowerdown => powerdn(3 DOWNTO 2),
		hipstatus => wire_receive_pcs1_hipstatus,
		invpol => wire_gnd,
		localrefclk => tx_localrefclk(1),
		masterclk => wire_gnd,
		parallelfdbk => wire_receive_pcs1_parallelfdbk,
		phfifordenable => rx_phfifordenable(1),
		phfifordenableout => wire_receive_pcs1_phfifordenableout,
		phfiforeset => rx_phfiforeset(1),
		phfiforesetout => wire_receive_pcs1_phfiforesetout,
		phfifowrdisable => rx_phfifowrdisable(1),
		phfifowrdisableout => wire_receive_pcs1_phfifowrdisableout,
		phfifox4bytesel => int_rx_phfifoxnbytesel(1),
		phfifox4rdenable => int_rx_phfifoxnrdenable(1),
		phfifox4wrclk => int_rx_phfifoxnwrclk(1),
		phfifox4wrenable => int_rx_phfifoxnwrenable(1),
		pipeenrevparallellpbkfromtx => int_pipeenrevparallellpbkfromtx(1),
		pipepowerdown => tx_pipepowerdownout(3 DOWNTO 2),
		pipepowerstate => tx_pipepowerstateout(7 DOWNTO 4),
		prbscidenable => rx_prbscidenable(1),
		quadreset => cent_unit_quadresetout(0),
		recoveredclk => rx_pma_clockout(1),
		refclk => refclk_pma(0),
		revbitorderwa => wire_gnd,
		revparallelfdbkdata => wire_receive_pcs1_revparallelfdbkdata,
		rmfifordena => wire_gnd,
		rmfiforeset => rx_rmfiforeset(1),
		rmfifowrena => wire_gnd,
		rxdetectvalid => tx_rxdetectvalidout(1),
		rxfound => rx_pcs_rxfound_wire(3 DOWNTO 2),
		signaldetected => rx_signaldetect_wire(1),
		xgmctrlin => wire_gnd,
		xgmdatain => wire_receive_pcs1_xgmdatain
	  );
	wire_receive_pcs2_hipelecidleinfersel <= (OTHERS => '0');
	wire_receive_pcs2_parallelfdbk <= (OTHERS => '0');
	wire_receive_pcs2_xgmdatain <= (OTHERS => '0');
	receive_pcs2 :  cycloneiv_hssi_rx_pcs
	  GENERIC MAP (
		align_pattern => "0101111100",
		align_pattern_length => 10,
		allow_align_polarity_inversion => "false",
		allow_pipe_polarity_inversion => "true",
		auto_spd_deassert_ph_fifo_rst_count => 8,
		auto_spd_phystatus_notify_count => 14,
		bit_slip_enable => "false",
		byte_order_invalid_code_or_run_disp_error => "true",
		byte_order_mode => "none",
		byte_order_pad_pattern => "0",
		byte_order_pattern => "0",
		byte_order_pld_ctrl_enable => "false",
		cdrctrl_bypass_ppm_detector_cycle => 1000,
		cdrctrl_cid_mode_enable => "true",
		cdrctrl_enable => "true",
		cdrctrl_mask_cycle => 800,
		cdrctrl_min_lock_to_ref_cycle => 63,
		cdrctrl_rxvalid_mask => "true",
		channel_bonding => "x4",
		channel_number => ((starting_channel_number + 2) MOD 4),
		channel_width => 8,
		clk1_mux_select => "recovered clock",
		clk2_mux_select => "digital reference clock",
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "pipe",
		dec_8b_10b_compatibility_mode => "true",
		dec_8b_10b_mode => "normal",
		deskew_pattern => "0",
		disable_auto_idle_insertion => "false",
		disable_running_disp_in_word_align => "false",
		disallow_kchar_after_pattern_ordered_set => "false",
		dprio_config_mode => "000001",
		elec_idle_gen1_sigdet_enable => "true",
		elec_idle_infer_enable => "false",
		elec_idle_num_com_detect => 3,
		enable_bit_reversal => "false",
		enable_self_test_mode => "false",
		force_signal_detect_dig => "true",
		hip_enable => "true",
		infiniband_invalid_code => 0,
		insert_pad_on_underflow => "false",
		num_align_code_groups_in_ordered_set => 0,
		num_align_cons_good_data => 16,
		num_align_cons_pat => 4,
		num_align_loss_sync_error => 17,
		ph_fifo_low_latency_enable => "true",
		ph_fifo_reg_mode => "true",
		protocol_hint => "pcie",
		rate_match_back_to_back => "false",
		rate_match_delete_threshold => 13,
		rate_match_empty_threshold => 5,
		rate_match_fifo_mode => "true",
		rate_match_full_threshold => 20,
		rate_match_insert_threshold => 11,
		rate_match_ordered_set_based => "false",
		rate_match_pattern1 => "11010000111010000011",
		rate_match_pattern2 => "00101111000101111100",
		rate_match_pattern_size => 20,
		rate_match_pipe_enable => "true",
		rate_match_reset_enable => "false",
		rate_match_skip_set_based => "true",
		rate_match_start_threshold => 7,
		rd_clk_mux_select => "int clock",
		recovered_clk_mux_select => "recovered clock",
		run_length => 40,
		run_length_enable => "true",
		rx_detect_bypass => "false",
		rx_phfifo_wait_cnt => 32,
		rxstatus_error_report_mode => 1,
		self_test_mode => "incremental",
		use_alignment_state_machine => "true",
		use_deskew_fifo => "false",
		use_double_data_mode => "false",
		use_parallel_loopback => "false"
	  )
	  PORT MAP ( 
		a1a2size => wire_gnd,
		alignstatus => wire_gnd,
		alignstatussync => wire_gnd,
		cdrctrlearlyeios => wire_receive_pcs2_cdrctrlearlyeios,
		cdrctrllocktorefclkout => wire_receive_pcs2_cdrctrllocktorefclkout,
		coreclkout => wire_receive_pcs2_coreclkout,
		datain => rx_pma_recoverdataout_wire(29 DOWNTO 20),
		digitalreset => rx_digitalreset_out(2),
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => rx_pcsdprioin_wire(1199 DOWNTO 800),
		dprioout => wire_receive_pcs2_dprioout,
		enabledeskew => wire_gnd,
		enabyteord => wire_gnd,
		enapatternalign => rx_enapatternalign(2),
		fifordin => wire_gnd,
		fiforesetrd => wire_gnd,
		hip8b10binvpolarity => pipe8b10binvpolarity(2),
		hipdataout => wire_receive_pcs2_hipdataout,
		hipdatavalid => wire_receive_pcs2_hipdatavalid,
		hipelecidle => wire_receive_pcs2_hipelecidle,
		hipelecidleinfersel => wire_receive_pcs2_hipelecidleinfersel,
		hipphydonestatus => wire_receive_pcs2_hipphydonestatus,
		hippowerdown => powerdn(5 DOWNTO 4),
		hipstatus => wire_receive_pcs2_hipstatus,
		invpol => wire_gnd,
		localrefclk => tx_localrefclk(2),
		masterclk => wire_gnd,
		parallelfdbk => wire_receive_pcs2_parallelfdbk,
		phfifordenable => rx_phfifordenable(2),
		phfifordenableout => wire_receive_pcs2_phfifordenableout,
		phfiforeset => rx_phfiforeset(2),
		phfiforesetout => wire_receive_pcs2_phfiforesetout,
		phfifowrdisable => rx_phfifowrdisable(2),
		phfifowrdisableout => wire_receive_pcs2_phfifowrdisableout,
		phfifox4bytesel => int_rx_phfifoxnbytesel(2),
		phfifox4rdenable => int_rx_phfifoxnrdenable(2),
		phfifox4wrclk => int_rx_phfifoxnwrclk(2),
		phfifox4wrenable => int_rx_phfifoxnwrenable(2),
		pipeenrevparallellpbkfromtx => int_pipeenrevparallellpbkfromtx(2),
		pipepowerdown => tx_pipepowerdownout(5 DOWNTO 4),
		pipepowerstate => tx_pipepowerstateout(11 DOWNTO 8),
		prbscidenable => rx_prbscidenable(2),
		quadreset => cent_unit_quadresetout(0),
		recoveredclk => rx_pma_clockout(2),
		refclk => refclk_pma(0),
		revbitorderwa => wire_gnd,
		revparallelfdbkdata => wire_receive_pcs2_revparallelfdbkdata,
		rmfifordena => wire_gnd,
		rmfiforeset => rx_rmfiforeset(2),
		rmfifowrena => wire_gnd,
		rxdetectvalid => tx_rxdetectvalidout(2),
		rxfound => rx_pcs_rxfound_wire(5 DOWNTO 4),
		signaldetected => rx_signaldetect_wire(2),
		xgmctrlin => wire_gnd,
		xgmdatain => wire_receive_pcs2_xgmdatain
	  );
	wire_receive_pcs3_hipelecidleinfersel <= (OTHERS => '0');
	wire_receive_pcs3_parallelfdbk <= (OTHERS => '0');
	wire_receive_pcs3_xgmdatain <= (OTHERS => '0');
	receive_pcs3 :  cycloneiv_hssi_rx_pcs
	  GENERIC MAP (
		align_pattern => "0101111100",
		align_pattern_length => 10,
		allow_align_polarity_inversion => "false",
		allow_pipe_polarity_inversion => "true",
		auto_spd_deassert_ph_fifo_rst_count => 8,
		auto_spd_phystatus_notify_count => 14,
		bit_slip_enable => "false",
		byte_order_invalid_code_or_run_disp_error => "true",
		byte_order_mode => "none",
		byte_order_pad_pattern => "0",
		byte_order_pattern => "0",
		byte_order_pld_ctrl_enable => "false",
		cdrctrl_bypass_ppm_detector_cycle => 1000,
		cdrctrl_cid_mode_enable => "true",
		cdrctrl_enable => "true",
		cdrctrl_mask_cycle => 800,
		cdrctrl_min_lock_to_ref_cycle => 63,
		cdrctrl_rxvalid_mask => "true",
		channel_bonding => "x4",
		channel_number => ((starting_channel_number + 3) MOD 4),
		channel_width => 8,
		clk1_mux_select => "recovered clock",
		clk2_mux_select => "digital reference clock",
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "pipe",
		dec_8b_10b_compatibility_mode => "true",
		dec_8b_10b_mode => "normal",
		deskew_pattern => "0",
		disable_auto_idle_insertion => "false",
		disable_running_disp_in_word_align => "false",
		disallow_kchar_after_pattern_ordered_set => "false",
		dprio_config_mode => "000001",
		elec_idle_gen1_sigdet_enable => "true",
		elec_idle_infer_enable => "false",
		elec_idle_num_com_detect => 3,
		enable_bit_reversal => "false",
		enable_self_test_mode => "false",
		force_signal_detect_dig => "true",
		hip_enable => "true",
		infiniband_invalid_code => 0,
		insert_pad_on_underflow => "false",
		num_align_code_groups_in_ordered_set => 0,
		num_align_cons_good_data => 16,
		num_align_cons_pat => 4,
		num_align_loss_sync_error => 17,
		ph_fifo_low_latency_enable => "true",
		ph_fifo_reg_mode => "true",
		protocol_hint => "pcie",
		rate_match_back_to_back => "false",
		rate_match_delete_threshold => 13,
		rate_match_empty_threshold => 5,
		rate_match_fifo_mode => "true",
		rate_match_full_threshold => 20,
		rate_match_insert_threshold => 11,
		rate_match_ordered_set_based => "false",
		rate_match_pattern1 => "11010000111010000011",
		rate_match_pattern2 => "00101111000101111100",
		rate_match_pattern_size => 20,
		rate_match_pipe_enable => "true",
		rate_match_reset_enable => "false",
		rate_match_skip_set_based => "true",
		rate_match_start_threshold => 7,
		rd_clk_mux_select => "int clock",
		recovered_clk_mux_select => "recovered clock",
		run_length => 40,
		run_length_enable => "true",
		rx_detect_bypass => "false",
		rx_phfifo_wait_cnt => 32,
		rxstatus_error_report_mode => 1,
		self_test_mode => "incremental",
		use_alignment_state_machine => "true",
		use_deskew_fifo => "false",
		use_double_data_mode => "false",
		use_parallel_loopback => "false"
	  )
	  PORT MAP ( 
		a1a2size => wire_gnd,
		alignstatus => wire_gnd,
		alignstatussync => wire_gnd,
		cdrctrlearlyeios => wire_receive_pcs3_cdrctrlearlyeios,
		cdrctrllocktorefclkout => wire_receive_pcs3_cdrctrllocktorefclkout,
		coreclkout => wire_receive_pcs3_coreclkout,
		datain => rx_pma_recoverdataout_wire(39 DOWNTO 30),
		digitalreset => rx_digitalreset_out(3),
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => rx_pcsdprioin_wire(1599 DOWNTO 1200),
		dprioout => wire_receive_pcs3_dprioout,
		enabledeskew => wire_gnd,
		enabyteord => wire_gnd,
		enapatternalign => rx_enapatternalign(3),
		fifordin => wire_gnd,
		fiforesetrd => wire_gnd,
		hip8b10binvpolarity => pipe8b10binvpolarity(3),
		hipdataout => wire_receive_pcs3_hipdataout,
		hipdatavalid => wire_receive_pcs3_hipdatavalid,
		hipelecidle => wire_receive_pcs3_hipelecidle,
		hipelecidleinfersel => wire_receive_pcs3_hipelecidleinfersel,
		hipphydonestatus => wire_receive_pcs3_hipphydonestatus,
		hippowerdown => powerdn(7 DOWNTO 6),
		hipstatus => wire_receive_pcs3_hipstatus,
		invpol => wire_gnd,
		localrefclk => tx_localrefclk(3),
		masterclk => wire_gnd,
		parallelfdbk => wire_receive_pcs3_parallelfdbk,
		phfifordenable => rx_phfifordenable(3),
		phfifordenableout => wire_receive_pcs3_phfifordenableout,
		phfiforeset => rx_phfiforeset(3),
		phfiforesetout => wire_receive_pcs3_phfiforesetout,
		phfifowrdisable => rx_phfifowrdisable(3),
		phfifowrdisableout => wire_receive_pcs3_phfifowrdisableout,
		phfifox4bytesel => int_rx_phfifoxnbytesel(3),
		phfifox4rdenable => int_rx_phfifoxnrdenable(3),
		phfifox4wrclk => int_rx_phfifoxnwrclk(3),
		phfifox4wrenable => int_rx_phfifoxnwrenable(3),
		pipeenrevparallellpbkfromtx => int_pipeenrevparallellpbkfromtx(3),
		pipepowerdown => tx_pipepowerdownout(7 DOWNTO 6),
		pipepowerstate => tx_pipepowerstateout(15 DOWNTO 12),
		prbscidenable => rx_prbscidenable(3),
		quadreset => cent_unit_quadresetout(0),
		recoveredclk => rx_pma_clockout(3),
		refclk => refclk_pma(0),
		revbitorderwa => wire_gnd,
		revparallelfdbkdata => wire_receive_pcs3_revparallelfdbkdata,
		rmfifordena => wire_gnd,
		rmfiforeset => rx_rmfiforeset(3),
		rmfifowrena => wire_gnd,
		rxdetectvalid => tx_rxdetectvalidout(3),
		rxfound => rx_pcs_rxfound_wire(7 DOWNTO 6),
		signaldetected => rx_signaldetect_wire(3),
		xgmctrlin => wire_gnd,
		xgmdatain => wire_receive_pcs3_xgmdatain
	  );
	wire_receive_pma0_w_lg_freqlocked613w(0) <= wire_receive_pma0_freqlocked AND wire_w_lg_w_rx_analogreset_range513w612w(0);
	wire_receive_pma0_locktodata <= wire_w_lg_w_lg_reconfig_togxb_busy514w601w(0);
	wire_w_lg_w_lg_reconfig_togxb_busy514w601w(0) <= wire_w_lg_reconfig_togxb_busy514w(0) AND rx_locktodata(0);
	wire_receive_pma0_testbussel <= "0110";
	receive_pma0 :  cycloneiv_hssi_rx_pma
	  GENERIC MAP (
		allow_serial_loopback => "false",
		channel_number => ((starting_channel_number + 0) MOD 4),
		common_mode => "0.82V",
		deserialization_factor => 10,
		dprio_config_mode => "000001",
		effective_data_rate => "2500 Mbps",
		enable_local_divider => "false",
		enable_ltd => "false",
		enable_ltr => "false",
		enable_second_order_loop => "false",
		eq_dc_gain => 3,
		eq_setting => 5,
		force_signal_detect => "false",
		logical_channel_address => (starting_channel_number + 0),
		loop_1_digital_filter => 8,
		offset_cancellation => 1,
		ppm_gen1_2_xcnt_en => 1,
		ppm_post_eidle => 0,
		ppmselect => 8,
		protocol_hint => "pcie",
		signal_detect_hysteresis => 4,
		signal_detect_hysteresis_valid_threshold => 14,
		signal_detect_loss_threshold => 3,
		termination => "OCT 100 Ohms",
		use_external_termination => "false"
	  )
	  PORT MAP ( 
		analogtestbus => wire_receive_pma0_analogtestbus,
		clockout => wire_receive_pma0_clockout,
		crupowerdn => cent_unit_rxcrupowerdn(0),
		datain => rx_datain(0),
		deserclock => rx_deserclock_in(0),
		diagnosticlpbkout => wire_receive_pma0_diagnosticlpbkout,
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => rx_pmadprioin_wire(299 DOWNTO 0),
		dprioout => wire_receive_pma0_dprioout,
		freqlocked => wire_receive_pma0_freqlocked,
		locktodata => wire_receive_pma0_locktodata,
		locktoref => rx_locktorefclk_wire(0),
		locktorefout => wire_receive_pma0_locktorefout,
		powerdn => cent_unit_rxibpowerdn(0),
		ppmdetectrefclk => rx_pll_pfdrefclkout_wire(0),
		recoverdataout => wire_receive_pma0_recoverdataout,
		reverselpbkout => wire_receive_pma0_reverselpbkout,
		rxpmareset => rx_analogreset_out(0),
		seriallpbkin => tx_serialloopbackout(0),
		signaldetect => wire_receive_pma0_signaldetect,
		testbussel => wire_receive_pma0_testbussel
	  );
	wire_receive_pma1_w_lg_freqlocked681w(0) <= wire_receive_pma1_freqlocked AND wire_w_lg_w_rx_analogreset_range513w612w(0);
	wire_receive_pma1_locktodata <= wire_w_lg_w_lg_reconfig_togxb_busy514w677w(0);
	wire_w_lg_w_lg_reconfig_togxb_busy514w677w(0) <= wire_w_lg_reconfig_togxb_busy514w(0) AND rx_locktodata(1);
	wire_receive_pma1_testbussel <= "0110";
	receive_pma1 :  cycloneiv_hssi_rx_pma
	  GENERIC MAP (
		allow_serial_loopback => "false",
		channel_number => ((starting_channel_number + 1) MOD 4),
		common_mode => "0.82V",
		deserialization_factor => 10,
		dprio_config_mode => "000001",
		effective_data_rate => "2500 Mbps",
		enable_local_divider => "false",
		enable_ltd => "false",
		enable_ltr => "false",
		enable_second_order_loop => "false",
		eq_dc_gain => 3,
		eq_setting => 5,
		force_signal_detect => "false",
		logical_channel_address => (starting_channel_number + 1),
		loop_1_digital_filter => 8,
		offset_cancellation => 1,
		ppm_gen1_2_xcnt_en => 1,
		ppm_post_eidle => 0,
		ppmselect => 8,
		protocol_hint => "pcie",
		signal_detect_hysteresis => 4,
		signal_detect_hysteresis_valid_threshold => 14,
		signal_detect_loss_threshold => 3,
		termination => "OCT 100 Ohms",
		use_external_termination => "false"
	  )
	  PORT MAP ( 
		analogtestbus => wire_receive_pma1_analogtestbus,
		clockout => wire_receive_pma1_clockout,
		crupowerdn => cent_unit_rxcrupowerdn(1),
		datain => rx_datain(1),
		deserclock => rx_deserclock_in(1),
		diagnosticlpbkout => wire_receive_pma1_diagnosticlpbkout,
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => rx_pmadprioin_wire(599 DOWNTO 300),
		dprioout => wire_receive_pma1_dprioout,
		freqlocked => wire_receive_pma1_freqlocked,
		locktodata => wire_receive_pma1_locktodata,
		locktoref => rx_locktorefclk_wire(1),
		locktorefout => wire_receive_pma1_locktorefout,
		powerdn => cent_unit_rxibpowerdn(1),
		ppmdetectrefclk => rx_pll_pfdrefclkout_wire(1),
		recoverdataout => wire_receive_pma1_recoverdataout,
		reverselpbkout => wire_receive_pma1_reverselpbkout,
		rxpmareset => rx_analogreset_out(1),
		seriallpbkin => tx_serialloopbackout(1),
		signaldetect => wire_receive_pma1_signaldetect,
		testbussel => wire_receive_pma1_testbussel
	  );
	wire_receive_pma2_w_lg_freqlocked748w(0) <= wire_receive_pma2_freqlocked AND wire_w_lg_w_rx_analogreset_range513w612w(0);
	wire_receive_pma2_locktodata <= wire_w_lg_w_lg_reconfig_togxb_busy514w744w(0);
	wire_w_lg_w_lg_reconfig_togxb_busy514w744w(0) <= wire_w_lg_reconfig_togxb_busy514w(0) AND rx_locktodata(2);
	wire_receive_pma2_testbussel <= "0110";
	receive_pma2 :  cycloneiv_hssi_rx_pma
	  GENERIC MAP (
		allow_serial_loopback => "false",
		channel_number => ((starting_channel_number + 2) MOD 4),
		common_mode => "0.82V",
		deserialization_factor => 10,
		dprio_config_mode => "000001",
		effective_data_rate => "2500 Mbps",
		enable_local_divider => "false",
		enable_ltd => "false",
		enable_ltr => "false",
		enable_second_order_loop => "false",
		eq_dc_gain => 3,
		eq_setting => 5,
		force_signal_detect => "false",
		logical_channel_address => (starting_channel_number + 2),
		loop_1_digital_filter => 8,
		offset_cancellation => 1,
		ppm_gen1_2_xcnt_en => 1,
		ppm_post_eidle => 0,
		ppmselect => 8,
		protocol_hint => "pcie",
		signal_detect_hysteresis => 4,
		signal_detect_hysteresis_valid_threshold => 14,
		signal_detect_loss_threshold => 3,
		termination => "OCT 100 Ohms",
		use_external_termination => "false"
	  )
	  PORT MAP ( 
		analogtestbus => wire_receive_pma2_analogtestbus,
		clockout => wire_receive_pma2_clockout,
		crupowerdn => cent_unit_rxcrupowerdn(2),
		datain => rx_datain(2),
		deserclock => rx_deserclock_in(2),
		diagnosticlpbkout => wire_receive_pma2_diagnosticlpbkout,
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => rx_pmadprioin_wire(899 DOWNTO 600),
		dprioout => wire_receive_pma2_dprioout,
		freqlocked => wire_receive_pma2_freqlocked,
		locktodata => wire_receive_pma2_locktodata,
		locktoref => rx_locktorefclk_wire(2),
		locktorefout => wire_receive_pma2_locktorefout,
		powerdn => cent_unit_rxibpowerdn(2),
		ppmdetectrefclk => rx_pll_pfdrefclkout_wire(2),
		recoverdataout => wire_receive_pma2_recoverdataout,
		reverselpbkout => wire_receive_pma2_reverselpbkout,
		rxpmareset => rx_analogreset_out(2),
		seriallpbkin => tx_serialloopbackout(2),
		signaldetect => wire_receive_pma2_signaldetect,
		testbussel => wire_receive_pma2_testbussel
	  );
	wire_receive_pma3_w_lg_freqlocked815w(0) <= wire_receive_pma3_freqlocked AND wire_w_lg_w_rx_analogreset_range513w612w(0);
	wire_receive_pma3_locktodata <= wire_w_lg_w_lg_reconfig_togxb_busy514w811w(0);
	wire_w_lg_w_lg_reconfig_togxb_busy514w811w(0) <= wire_w_lg_reconfig_togxb_busy514w(0) AND rx_locktodata(3);
	wire_receive_pma3_testbussel <= "0110";
	receive_pma3 :  cycloneiv_hssi_rx_pma
	  GENERIC MAP (
		allow_serial_loopback => "false",
		channel_number => ((starting_channel_number + 3) MOD 4),
		common_mode => "0.82V",
		deserialization_factor => 10,
		dprio_config_mode => "000001",
		effective_data_rate => "2500 Mbps",
		enable_local_divider => "false",
		enable_ltd => "false",
		enable_ltr => "false",
		enable_second_order_loop => "false",
		eq_dc_gain => 3,
		eq_setting => 5,
		force_signal_detect => "false",
		logical_channel_address => (starting_channel_number + 3),
		loop_1_digital_filter => 8,
		offset_cancellation => 1,
		ppm_gen1_2_xcnt_en => 1,
		ppm_post_eidle => 0,
		ppmselect => 8,
		protocol_hint => "pcie",
		signal_detect_hysteresis => 4,
		signal_detect_hysteresis_valid_threshold => 14,
		signal_detect_loss_threshold => 3,
		termination => "OCT 100 Ohms",
		use_external_termination => "false"
	  )
	  PORT MAP ( 
		analogtestbus => wire_receive_pma3_analogtestbus,
		clockout => wire_receive_pma3_clockout,
		crupowerdn => cent_unit_rxcrupowerdn(3),
		datain => rx_datain(3),
		deserclock => rx_deserclock_in(3),
		diagnosticlpbkout => wire_receive_pma3_diagnosticlpbkout,
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => rx_pmadprioin_wire(1199 DOWNTO 900),
		dprioout => wire_receive_pma3_dprioout,
		freqlocked => wire_receive_pma3_freqlocked,
		locktodata => wire_receive_pma3_locktodata,
		locktoref => rx_locktorefclk_wire(3),
		locktorefout => wire_receive_pma3_locktorefout,
		powerdn => cent_unit_rxibpowerdn(3),
		ppmdetectrefclk => rx_pll_pfdrefclkout_wire(3),
		recoverdataout => wire_receive_pma3_recoverdataout,
		reverselpbkout => wire_receive_pma3_reverselpbkout,
		rxpmareset => rx_analogreset_out(3),
		seriallpbkin => tx_serialloopbackout(3),
		signaldetect => wire_receive_pma3_signaldetect,
		testbussel => wire_receive_pma3_testbussel
	  );
	wire_transmit_pcs0_ctrlenable <= ( "0" & "0");
	wire_transmit_pcs0_datainfull <= (OTHERS => '0');
	wire_transmit_pcs0_dispval <= ( "0" & "0");
	wire_transmit_pcs0_forcedisp <= ( "0" & "0");
	wire_transmit_pcs0_hipdatain <= ( tx_forcedispcompliance(0) & tx_ctrlenable(0) & tx_datain_wire(7 DOWNTO 0));
	transmit_pcs0 :  cycloneiv_hssi_tx_pcs
	  GENERIC MAP (
		allow_polarity_inversion => "false",
		bitslip_enable => "false",
		channel_bonding => "x4",
		channel_number => ((starting_channel_number + 0) MOD 4),
		channel_width => 8,
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "pipe",
		disable_ph_low_latency_mode => "false",
		disparity_mode => "new",
		dprio_config_mode => "000001",
		elec_idle_delay => 4,
		enable_bit_reversal => "false",
		enable_idle_selection => "false",
		enable_reverse_parallel_loopback => "true",
		enable_self_test_mode => "false",
		enc_8b_10b_compatibility_mode => "true",
		enc_8b_10b_mode => "normal",
		hip_enable => "true",
		ph_fifo_reg_mode => "true",
		prbs_cid_pattern => "false",
		protocol_hint => "pcie",
		refclk_select => "central",
		self_test_mode => "incremental",
		use_double_data_mode => "false",
		wr_clk_mux_select => "int_clk"
	  )
	  PORT MAP ( 
		coreclkout => wire_transmit_pcs0_coreclkout,
		ctrlenable => wire_transmit_pcs0_ctrlenable,
		datainfull => wire_transmit_pcs0_datainfull,
		dataout => wire_transmit_pcs0_dataout,
		digitalreset => tx_digitalreset_out(0),
		dispval => wire_transmit_pcs0_dispval,
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => tx_dprioin_wire(149 DOWNTO 0),
		dprioout => wire_transmit_pcs0_dprioout,
		enrevparallellpbk => tx_revparallellpbken(0),
		forcedisp => wire_transmit_pcs0_forcedisp,
		forceelecidleout => wire_transmit_pcs0_forceelecidleout,
		grayelecidleinferselout => wire_transmit_pcs0_grayelecidleinferselout,
		hipdatain => wire_transmit_pcs0_hipdatain,
		hipdetectrxloop => tx_detectrxloop(0),
		hipelecidleinfersel => rx_elecidleinfersel(2 DOWNTO 0),
		hipforceelecidle => tx_forceelecidle(0),
		hippowerdn => powerdn(1 DOWNTO 0),
		invpol => tx_invpolarity(0),
		localrefclk => tx_localrefclk(0),
		phfiforddisable => wire_gnd,
		phfiforddisableout => wire_transmit_pcs0_phfiforddisableout,
		phfiforeset => tx_phfiforeset(0),
		phfiforesetout => wire_transmit_pcs0_phfiforesetout,
		phfifowrenable => wire_vcc,
		phfifowrenableout => wire_transmit_pcs0_phfifowrenableout,
		phfifox4bytesel => int_tx_phfifoxnbytesel(0),
		phfifox4rdclk => int_tx_phfifoxnrdclk(0),
		phfifox4rdenable => int_tx_phfifoxnrdenable(0),
		phfifox4wrenable => int_tx_phfifoxnwrenable(0),
		pipeenrevparallellpbkout => wire_transmit_pcs0_pipeenrevparallellpbkout,
		pipepowerdownout => wire_transmit_pcs0_pipepowerdownout,
		pipepowerstateout => wire_transmit_pcs0_pipepowerstateout,
		pipestatetransdone => wire_gnd,
		quadreset => cent_unit_quadresetout(0),
		refclk => refclk_pma(0),
		revparallelfdbk => rx_revparallelfdbkdata(19 DOWNTO 0),
		txdetectrx => wire_transmit_pcs0_txdetectrx
	  );
	wire_transmit_pcs1_ctrlenable <= ( "0" & "0");
	wire_transmit_pcs1_datainfull <= (OTHERS => '0');
	wire_transmit_pcs1_dispval <= ( "0" & "0");
	wire_transmit_pcs1_forcedisp <= ( "0" & "0");
	wire_transmit_pcs1_hipdatain <= ( tx_forcedispcompliance(1) & tx_ctrlenable(1) & tx_datain_wire(15 DOWNTO 8));
	transmit_pcs1 :  cycloneiv_hssi_tx_pcs
	  GENERIC MAP (
		allow_polarity_inversion => "false",
		bitslip_enable => "false",
		channel_bonding => "x4",
		channel_number => ((starting_channel_number + 1) MOD 4),
		channel_width => 8,
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "pipe",
		disable_ph_low_latency_mode => "false",
		disparity_mode => "new",
		dprio_config_mode => "000001",
		elec_idle_delay => 4,
		enable_bit_reversal => "false",
		enable_idle_selection => "false",
		enable_reverse_parallel_loopback => "true",
		enable_self_test_mode => "false",
		enc_8b_10b_compatibility_mode => "true",
		enc_8b_10b_mode => "normal",
		hip_enable => "true",
		ph_fifo_reg_mode => "true",
		prbs_cid_pattern => "false",
		protocol_hint => "pcie",
		refclk_select => "central",
		self_test_mode => "incremental",
		use_double_data_mode => "false",
		wr_clk_mux_select => "int_clk"
	  )
	  PORT MAP ( 
		coreclkout => wire_transmit_pcs1_coreclkout,
		ctrlenable => wire_transmit_pcs1_ctrlenable,
		datainfull => wire_transmit_pcs1_datainfull,
		dataout => wire_transmit_pcs1_dataout,
		digitalreset => tx_digitalreset_out(1),
		dispval => wire_transmit_pcs1_dispval,
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => tx_dprioin_wire(299 DOWNTO 150),
		dprioout => wire_transmit_pcs1_dprioout,
		enrevparallellpbk => tx_revparallellpbken(1),
		forcedisp => wire_transmit_pcs1_forcedisp,
		forceelecidleout => wire_transmit_pcs1_forceelecidleout,
		grayelecidleinferselout => wire_transmit_pcs1_grayelecidleinferselout,
		hipdatain => wire_transmit_pcs1_hipdatain,
		hipdetectrxloop => tx_detectrxloop(1),
		hipelecidleinfersel => rx_elecidleinfersel(5 DOWNTO 3),
		hipforceelecidle => tx_forceelecidle(1),
		hippowerdn => powerdn(3 DOWNTO 2),
		invpol => tx_invpolarity(1),
		localrefclk => tx_localrefclk(1),
		phfiforddisable => wire_gnd,
		phfiforddisableout => wire_transmit_pcs1_phfiforddisableout,
		phfiforeset => tx_phfiforeset(1),
		phfiforesetout => wire_transmit_pcs1_phfiforesetout,
		phfifowrenable => wire_vcc,
		phfifowrenableout => wire_transmit_pcs1_phfifowrenableout,
		phfifox4bytesel => int_tx_phfifoxnbytesel(1),
		phfifox4rdclk => int_tx_phfifoxnrdclk(1),
		phfifox4rdenable => int_tx_phfifoxnrdenable(1),
		phfifox4wrenable => int_tx_phfifoxnwrenable(1),
		pipeenrevparallellpbkout => wire_transmit_pcs1_pipeenrevparallellpbkout,
		pipepowerdownout => wire_transmit_pcs1_pipepowerdownout,
		pipepowerstateout => wire_transmit_pcs1_pipepowerstateout,
		pipestatetransdone => wire_gnd,
		quadreset => cent_unit_quadresetout(0),
		refclk => refclk_pma(0),
		revparallelfdbk => rx_revparallelfdbkdata(39 DOWNTO 20),
		txdetectrx => wire_transmit_pcs1_txdetectrx
	  );
	wire_transmit_pcs2_ctrlenable <= ( "0" & "0");
	wire_transmit_pcs2_datainfull <= (OTHERS => '0');
	wire_transmit_pcs2_dispval <= ( "0" & "0");
	wire_transmit_pcs2_forcedisp <= ( "0" & "0");
	wire_transmit_pcs2_hipdatain <= ( tx_forcedispcompliance(2) & tx_ctrlenable(2) & tx_datain_wire(23 DOWNTO 16));
	transmit_pcs2 :  cycloneiv_hssi_tx_pcs
	  GENERIC MAP (
		allow_polarity_inversion => "false",
		bitslip_enable => "false",
		channel_bonding => "x4",
		channel_number => ((starting_channel_number + 2) MOD 4),
		channel_width => 8,
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "pipe",
		disable_ph_low_latency_mode => "false",
		disparity_mode => "new",
		dprio_config_mode => "000001",
		elec_idle_delay => 4,
		enable_bit_reversal => "false",
		enable_idle_selection => "false",
		enable_reverse_parallel_loopback => "true",
		enable_self_test_mode => "false",
		enc_8b_10b_compatibility_mode => "true",
		enc_8b_10b_mode => "normal",
		hip_enable => "true",
		ph_fifo_reg_mode => "true",
		prbs_cid_pattern => "false",
		protocol_hint => "pcie",
		refclk_select => "central",
		self_test_mode => "incremental",
		use_double_data_mode => "false",
		wr_clk_mux_select => "int_clk"
	  )
	  PORT MAP ( 
		coreclkout => wire_transmit_pcs2_coreclkout,
		ctrlenable => wire_transmit_pcs2_ctrlenable,
		datainfull => wire_transmit_pcs2_datainfull,
		dataout => wire_transmit_pcs2_dataout,
		digitalreset => tx_digitalreset_out(2),
		dispval => wire_transmit_pcs2_dispval,
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => tx_dprioin_wire(449 DOWNTO 300),
		dprioout => wire_transmit_pcs2_dprioout,
		enrevparallellpbk => tx_revparallellpbken(2),
		forcedisp => wire_transmit_pcs2_forcedisp,
		forceelecidleout => wire_transmit_pcs2_forceelecidleout,
		grayelecidleinferselout => wire_transmit_pcs2_grayelecidleinferselout,
		hipdatain => wire_transmit_pcs2_hipdatain,
		hipdetectrxloop => tx_detectrxloop(2),
		hipelecidleinfersel => rx_elecidleinfersel(8 DOWNTO 6),
		hipforceelecidle => tx_forceelecidle(2),
		hippowerdn => powerdn(5 DOWNTO 4),
		invpol => tx_invpolarity(2),
		localrefclk => tx_localrefclk(2),
		phfiforddisable => wire_gnd,
		phfiforddisableout => wire_transmit_pcs2_phfiforddisableout,
		phfiforeset => tx_phfiforeset(2),
		phfiforesetout => wire_transmit_pcs2_phfiforesetout,
		phfifowrenable => wire_vcc,
		phfifowrenableout => wire_transmit_pcs2_phfifowrenableout,
		phfifox4bytesel => int_tx_phfifoxnbytesel(2),
		phfifox4rdclk => int_tx_phfifoxnrdclk(2),
		phfifox4rdenable => int_tx_phfifoxnrdenable(2),
		phfifox4wrenable => int_tx_phfifoxnwrenable(2),
		pipeenrevparallellpbkout => wire_transmit_pcs2_pipeenrevparallellpbkout,
		pipepowerdownout => wire_transmit_pcs2_pipepowerdownout,
		pipepowerstateout => wire_transmit_pcs2_pipepowerstateout,
		pipestatetransdone => wire_gnd,
		quadreset => cent_unit_quadresetout(0),
		refclk => refclk_pma(0),
		revparallelfdbk => rx_revparallelfdbkdata(59 DOWNTO 40),
		txdetectrx => wire_transmit_pcs2_txdetectrx
	  );
	wire_transmit_pcs3_ctrlenable <= ( "0" & "0");
	wire_transmit_pcs3_datainfull <= (OTHERS => '0');
	wire_transmit_pcs3_dispval <= ( "0" & "0");
	wire_transmit_pcs3_forcedisp <= ( "0" & "0");
	wire_transmit_pcs3_hipdatain <= ( tx_forcedispcompliance(3) & tx_ctrlenable(3) & tx_datain_wire(31 DOWNTO 24));
	transmit_pcs3 :  cycloneiv_hssi_tx_pcs
	  GENERIC MAP (
		allow_polarity_inversion => "false",
		bitslip_enable => "false",
		channel_bonding => "x4",
		channel_number => ((starting_channel_number + 3) MOD 4),
		channel_width => 8,
		core_clock_0ppm => "false",
		datapath_low_latency_mode => "false",
		datapath_protocol => "pipe",
		disable_ph_low_latency_mode => "false",
		disparity_mode => "new",
		dprio_config_mode => "000001",
		elec_idle_delay => 4,
		enable_bit_reversal => "false",
		enable_idle_selection => "false",
		enable_reverse_parallel_loopback => "true",
		enable_self_test_mode => "false",
		enc_8b_10b_compatibility_mode => "true",
		enc_8b_10b_mode => "normal",
		hip_enable => "true",
		ph_fifo_reg_mode => "true",
		prbs_cid_pattern => "false",
		protocol_hint => "pcie",
		refclk_select => "central",
		self_test_mode => "incremental",
		use_double_data_mode => "false",
		wr_clk_mux_select => "int_clk"
	  )
	  PORT MAP ( 
		coreclkout => wire_transmit_pcs3_coreclkout,
		ctrlenable => wire_transmit_pcs3_ctrlenable,
		datainfull => wire_transmit_pcs3_datainfull,
		dataout => wire_transmit_pcs3_dataout,
		digitalreset => tx_digitalreset_out(3),
		dispval => wire_transmit_pcs3_dispval,
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => tx_dprioin_wire(599 DOWNTO 450),
		dprioout => wire_transmit_pcs3_dprioout,
		enrevparallellpbk => tx_revparallellpbken(3),
		forcedisp => wire_transmit_pcs3_forcedisp,
		forceelecidleout => wire_transmit_pcs3_forceelecidleout,
		grayelecidleinferselout => wire_transmit_pcs3_grayelecidleinferselout,
		hipdatain => wire_transmit_pcs3_hipdatain,
		hipdetectrxloop => tx_detectrxloop(3),
		hipelecidleinfersel => rx_elecidleinfersel(11 DOWNTO 9),
		hipforceelecidle => tx_forceelecidle(3),
		hippowerdn => powerdn(7 DOWNTO 6),
		invpol => tx_invpolarity(3),
		localrefclk => tx_localrefclk(3),
		phfiforddisable => wire_gnd,
		phfiforddisableout => wire_transmit_pcs3_phfiforddisableout,
		phfiforeset => tx_phfiforeset(3),
		phfiforesetout => wire_transmit_pcs3_phfiforesetout,
		phfifowrenable => wire_vcc,
		phfifowrenableout => wire_transmit_pcs3_phfifowrenableout,
		phfifox4bytesel => int_tx_phfifoxnbytesel(3),
		phfifox4rdclk => int_tx_phfifoxnrdclk(3),
		phfifox4rdenable => int_tx_phfifoxnrdenable(3),
		phfifox4wrenable => int_tx_phfifoxnwrenable(3),
		pipeenrevparallellpbkout => wire_transmit_pcs3_pipeenrevparallellpbkout,
		pipepowerdownout => wire_transmit_pcs3_pipepowerdownout,
		pipepowerstateout => wire_transmit_pcs3_pipepowerstateout,
		pipestatetransdone => wire_gnd,
		quadreset => cent_unit_quadresetout(0),
		refclk => refclk_pma(0),
		revparallelfdbk => rx_revparallelfdbkdata(79 DOWNTO 60),
		txdetectrx => wire_transmit_pcs3_txdetectrx
	  );
	wire_transmit_pma0_datain <= ( tx_dataout_pcs_to_pma(9 DOWNTO 0));
	transmit_pma0 :  cycloneiv_hssi_tx_pma
	  GENERIC MAP (
		channel_number => ((starting_channel_number + 0) MOD 4),
		common_mode => "0.65V",
		dprio_config_mode => "000001",
		effective_data_rate => "2500 Mbps",
		enable_diagnostic_loopback => "false",
		enable_reverse_serial_loopback => "false",
		logical_channel_address => (starting_channel_number + 0),
		preemp_tap_1 => 1,
		protocol_hint => "pcie",
		rx_detect => 0,
		serialization_factor => 10,
		slew_rate => "low",
		termination => "OCT 100 Ohms",
		use_external_termination => "false",
		use_rx_detect => "true",
		vod_selection => 4
	  )
	  PORT MAP ( 
		cgbpowerdn => cent_unit_txdividerpowerdown(0),
		clockout => wire_transmit_pma0_clockout,
		datain => wire_transmit_pma0_datain,
		dataout => wire_transmit_pma0_dataout,
		detectrxpowerdown => cent_unit_txdetectrxpowerdn(0),
		diagnosticlpbkin => tx_diagnosticlpbkin(0),
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => tx_pmadprioin_wire(299 DOWNTO 0),
		dprioout => wire_transmit_pma0_dprioout,
		fastrefclk0in => tx_pma_fastrefclk0in(0),
		forceelecidle => tx_pcs_forceelecidleout(0),
		powerdn => cent_unit_txobpowerdn(0),
		refclk0in => tx_pma_refclk0in(0),
		refclk0inpulse => tx_pma_refclk0inpulse(0),
		reverselpbkin => rx_reverselpbkout(0),
		rxdetecten => txdetectrxout(0),
		rxdetectvalidout => wire_transmit_pma0_rxdetectvalidout,
		rxfoundout => wire_transmit_pma0_rxfoundout,
		seriallpbkout => wire_transmit_pma0_seriallpbkout,
		txpmareset => tx_analogreset_out(0)
	  );
	wire_transmit_pma1_datain <= ( tx_dataout_pcs_to_pma(19 DOWNTO 10));
	transmit_pma1 :  cycloneiv_hssi_tx_pma
	  GENERIC MAP (
		channel_number => ((starting_channel_number + 1) MOD 4),
		common_mode => "0.65V",
		dprio_config_mode => "000001",
		effective_data_rate => "2500 Mbps",
		enable_diagnostic_loopback => "false",
		enable_reverse_serial_loopback => "false",
		logical_channel_address => (starting_channel_number + 1),
		preemp_tap_1 => 1,
		protocol_hint => "pcie",
		rx_detect => 0,
		serialization_factor => 10,
		slew_rate => "low",
		termination => "OCT 100 Ohms",
		use_external_termination => "false",
		use_rx_detect => "true",
		vod_selection => 4
	  )
	  PORT MAP ( 
		cgbpowerdn => cent_unit_txdividerpowerdown(1),
		clockout => wire_transmit_pma1_clockout,
		datain => wire_transmit_pma1_datain,
		dataout => wire_transmit_pma1_dataout,
		detectrxpowerdown => cent_unit_txdetectrxpowerdn(1),
		diagnosticlpbkin => tx_diagnosticlpbkin(1),
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => tx_pmadprioin_wire(599 DOWNTO 300),
		dprioout => wire_transmit_pma1_dprioout,
		fastrefclk0in => tx_pma_fastrefclk0in(1),
		forceelecidle => tx_pcs_forceelecidleout(1),
		powerdn => cent_unit_txobpowerdn(1),
		refclk0in => tx_pma_refclk0in(1),
		refclk0inpulse => tx_pma_refclk0inpulse(1),
		reverselpbkin => rx_reverselpbkout(1),
		rxdetecten => txdetectrxout(1),
		rxdetectvalidout => wire_transmit_pma1_rxdetectvalidout,
		rxfoundout => wire_transmit_pma1_rxfoundout,
		seriallpbkout => wire_transmit_pma1_seriallpbkout,
		txpmareset => tx_analogreset_out(1)
	  );
	wire_transmit_pma2_datain <= ( tx_dataout_pcs_to_pma(29 DOWNTO 20));
	transmit_pma2 :  cycloneiv_hssi_tx_pma
	  GENERIC MAP (
		channel_number => ((starting_channel_number + 2) MOD 4),
		common_mode => "0.65V",
		dprio_config_mode => "000001",
		effective_data_rate => "2500 Mbps",
		enable_diagnostic_loopback => "false",
		enable_reverse_serial_loopback => "false",
		logical_channel_address => (starting_channel_number + 2),
		preemp_tap_1 => 1,
		protocol_hint => "pcie",
		rx_detect => 0,
		serialization_factor => 10,
		slew_rate => "low",
		termination => "OCT 100 Ohms",
		use_external_termination => "false",
		use_rx_detect => "true",
		vod_selection => 4
	  )
	  PORT MAP ( 
		cgbpowerdn => cent_unit_txdividerpowerdown(2),
		clockout => wire_transmit_pma2_clockout,
		datain => wire_transmit_pma2_datain,
		dataout => wire_transmit_pma2_dataout,
		detectrxpowerdown => cent_unit_txdetectrxpowerdn(2),
		diagnosticlpbkin => tx_diagnosticlpbkin(2),
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => tx_pmadprioin_wire(899 DOWNTO 600),
		dprioout => wire_transmit_pma2_dprioout,
		fastrefclk0in => tx_pma_fastrefclk0in(2),
		forceelecidle => tx_pcs_forceelecidleout(2),
		powerdn => cent_unit_txobpowerdn(2),
		refclk0in => tx_pma_refclk0in(2),
		refclk0inpulse => tx_pma_refclk0inpulse(2),
		reverselpbkin => rx_reverselpbkout(2),
		rxdetecten => txdetectrxout(2),
		rxdetectvalidout => wire_transmit_pma2_rxdetectvalidout,
		rxfoundout => wire_transmit_pma2_rxfoundout,
		seriallpbkout => wire_transmit_pma2_seriallpbkout,
		txpmareset => tx_analogreset_out(2)
	  );
	wire_transmit_pma3_datain <= ( tx_dataout_pcs_to_pma(39 DOWNTO 30));
	transmit_pma3 :  cycloneiv_hssi_tx_pma
	  GENERIC MAP (
		channel_number => ((starting_channel_number + 3) MOD 4),
		common_mode => "0.65V",
		dprio_config_mode => "000001",
		effective_data_rate => "2500 Mbps",
		enable_diagnostic_loopback => "false",
		enable_reverse_serial_loopback => "false",
		logical_channel_address => (starting_channel_number + 3),
		preemp_tap_1 => 1,
		protocol_hint => "pcie",
		rx_detect => 0,
		serialization_factor => 10,
		slew_rate => "low",
		termination => "OCT 100 Ohms",
		use_external_termination => "false",
		use_rx_detect => "true",
		vod_selection => 4
	  )
	  PORT MAP ( 
		cgbpowerdn => cent_unit_txdividerpowerdown(3),
		clockout => wire_transmit_pma3_clockout,
		datain => wire_transmit_pma3_datain,
		dataout => wire_transmit_pma3_dataout,
		detectrxpowerdown => cent_unit_txdetectrxpowerdn(3),
		diagnosticlpbkin => tx_diagnosticlpbkin(3),
		dpriodisable => w_cent_unit_dpriodisableout1w(0),
		dprioin => tx_pmadprioin_wire(1199 DOWNTO 900),
		dprioout => wire_transmit_pma3_dprioout,
		fastrefclk0in => tx_pma_fastrefclk0in(3),
		forceelecidle => tx_pcs_forceelecidleout(3),
		powerdn => cent_unit_txobpowerdn(3),
		refclk0in => tx_pma_refclk0in(3),
		refclk0inpulse => tx_pma_refclk0inpulse(3),
		reverselpbkin => rx_reverselpbkout(3),
		rxdetecten => txdetectrxout(3),
		rxdetectvalidout => wire_transmit_pma3_rxdetectvalidout,
		rxfoundout => wire_transmit_pma3_rxfoundout,
		seriallpbkout => wire_transmit_pma3_seriallpbkout,
		txpmareset => tx_analogreset_out(3)
	  );
	PROCESS (fixedclk)
	BEGIN
		IF (fixedclk = '1' AND fixedclk'event) THEN fixedclk_div <= (NOT fixedclk_div_in);
		END IF;
	END PROCESS;
	PROCESS (fixedclk)
	BEGIN
		IF (fixedclk = '0' AND fixedclk'event) THEN reconfig_togxb_busy_reg <= ( reconfig_togxb_busy_reg(0) & reconfig_togxb_busy);
		END IF;
	END PROCESS;

 END RTL; --Hard_IP_x4_serdes_alt_c3gxb_41f8
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Hard_IP_x4_serdes IS
	GENERIC
	(
		starting_channel_number		: NATURAL := 0
	);
	PORT
	(
		cal_blk_clk		: IN STD_LOGIC ;
		fixedclk		: IN STD_LOGIC ;
		gxb_powerdown		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		pipe8b10binvpolarity		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		pll_areset		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		pll_inclk		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		powerdn		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		reconfig_clk		: IN STD_LOGIC ;
		reconfig_togxb		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		rx_analogreset		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		rx_datain		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		rx_digitalreset		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		rx_elecidleinfersel		: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
		tx_ctrlenable		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		tx_datain		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		tx_detectrxloop		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		tx_digitalreset		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		tx_forcedispcompliance		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		tx_forceelecidle		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		coreclkout		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		hip_tx_clkout		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		pipedatavalid		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		pipeelecidle		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		pipephydonestatus		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		pipestatus		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
		pll_locked		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		reconfig_fromgxb		: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
		rx_ctrldetect		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		rx_dataout		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
		rx_freqlocked		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		rx_patterndetect		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		rx_syncstatus		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		tx_dataout		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
END Hard_IP_x4_serdes;


ARCHITECTURE RTL OF hard_ip_x4_serdes IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "alt_c3gxb";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "effective_data_rate=2500 Mbps;enable_lc_tx_pll=false;enable_pll_inclk_alt_drive_rx_cru=true;enable_pll_inclk_drive_rx_cru=true;equalizer_dcgain_setting=1;gen_reconfig_pll=false;gx_channel_type=;input_clock_frequency=100.0 MHz;intended_device_family=Cyclone IV GX;intended_device_speed_grade=6;intended_device_variant=ANY;loopback_mode=none;lpm_type=alt_c3gxb;number_of_channels=4;operation_mode=duplex;pll_bandwidth_type=Auto;pll_control_width=1;pll_inclk_period=10000;pll_pfd_fb_mode=internal;preemphasis_ctrl_1stposttap_setting=1;protocol=pcie;receiver_termination=oct_100_ohms;reconfig_dprio_mode=0;rx_8b_10b_mode=normal;rx_align_pattern=0101111100;rx_align_pattern_length=10;rx_allow_align_polarity_inversion=false;rx_allow_pipe_polarity_inversion=true;rx_bitslip_enable=false;rx_byte_ordering_mode=NONE;rx_channel_bonding=x4;rx_channel_width=8;rx_common_mode=0.82v;rx_cru_inclock0_period=10000;rx_datapath_protocol=pipe;rx_data_rate=2500;rx_data_rate_remainder=0;rx_digitalreset_port_width=1;rx_enable_bit_reversal=false;rx_enable_lock_to_data_sig=false;rx_enable_lock_to_refclk_sig=false;rx_enable_self_test_mode=false;rx_force_signal_detect=false;rx_ppmselect=8;rx_rate_match_fifo_mode=normal;rx_rate_match_pattern1=11010000111010000011;rx_rate_match_pattern2=00101111000101111100;rx_rate_match_pattern_size=20;rx_run_length=40;rx_run_length_enable=true;rx_signal_detect_threshold=4;rx_use_align_state_machine=true;rx_use_clkout=false;rx_use_coreclk=false;" & 
	                                                    "rx_use_deserializer_double_data_mode=false;rx_use_deskew_fifo=false;rx_use_double_data_mode=false;rx_use_pipe8b10binvpolarity=true;rx_use_rate_match_pattern1_only=false;transmitter_termination=oct_100_ohms;tx_8b_10b_mode=normal;tx_allow_polarity_inversion=false;tx_channel_bonding=x4;tx_channel_width=8;tx_clkout_width=4;tx_common_mode=0.65v;tx_data_rate=2500;tx_data_rate_remainder=0;tx_digitalreset_port_width=1;tx_enable_bit_reversal=false;tx_enable_self_test_mode=false;tx_pll_bandwidth_type=Auto;tx_pll_inclk0_period=10000;tx_pll_type=CMU;tx_slew_rate=low;tx_transmit_protocol=pipe;tx_use_coreclk=false;tx_use_double_data_mode=false;tx_use_serializer_double_data_mode=false;use_calibration_block=true;vod_ctrl_setting=4;coreclkout_control_width=1;elec_idle_infer_enable=false;enable_0ppm=false;equalization_setting=5;gxb_powerdown_width=1;hip_enable=true;iqtxrxclk_allowed=;number_of_quads=1;pll_divide_by=2;pll_multiply_by=25;reconfig_calibration=true;reconfig_fromgxb_port_width=5;reconfig_pll_control_width=1;reconfig_togxb_port_width=4;rx_cdrctrl_enable=true;rx_deskew_pattern=0;rx_dwidth_factor=1;rx_enable_second_order_loop=false;rx_loop_1_digital_filter=8;rx_signal_detect_loss_threshold=3;rx_signal_detect_valid_threshold=14;rx_use_external_termination=false;rx_word_aligner_num_byte=1;top_module_name=Hard_IP_x4_serdes;tx_bitslip_enable=FALSE;tx_dwidth_factor=1;tx_use_external_termination=false;";
	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (11 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (4 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire12	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire13	: STD_LOGIC_VECTOR (3 DOWNTO 0);



	COMPONENT Hard_IP_x4_serdes_alt_c3gxb_41f8
	GENERIC (
		starting_channel_number		: NATURAL
	);
	PORT (
			cal_blk_clk	: IN STD_LOGIC ;
			fixedclk	: IN STD_LOGIC ;
			gxb_powerdown	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			pipe8b10binvpolarity	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			pll_areset	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			pll_inclk	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			powerdn	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			reconfig_clk	: IN STD_LOGIC ;
			reconfig_togxb	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			rx_analogreset	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_datain	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			rx_digitalreset	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			rx_elecidleinfersel	: IN STD_LOGIC_VECTOR (11 DOWNTO 0);
			tx_ctrlenable	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			tx_datain	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			tx_detectrxloop	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			tx_digitalreset	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			tx_forcedispcompliance	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			tx_forceelecidle	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			coreclkout	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			hip_tx_clkout	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			pipedatavalid	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			pipeelecidle	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			pipephydonestatus	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			pipestatus	: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
			pll_locked	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			reconfig_fromgxb	: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
			rx_ctrldetect	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			rx_dataout	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			rx_freqlocked	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			rx_patterndetect	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			rx_syncstatus	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			tx_dataout	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	coreclkout    <= sub_wire0(0 DOWNTO 0);
	hip_tx_clkout    <= sub_wire1(3 DOWNTO 0);
	pipedatavalid    <= sub_wire2(3 DOWNTO 0);
	pipeelecidle    <= sub_wire3(3 DOWNTO 0);
	pipephydonestatus    <= sub_wire4(3 DOWNTO 0);
	pipestatus    <= sub_wire5(11 DOWNTO 0);
	pll_locked    <= sub_wire6(0 DOWNTO 0);
	reconfig_fromgxb    <= sub_wire7(4 DOWNTO 0);
	rx_ctrldetect    <= sub_wire8(3 DOWNTO 0);
	rx_dataout    <= sub_wire9(31 DOWNTO 0);
	rx_freqlocked    <= sub_wire10(3 DOWNTO 0);
	rx_patterndetect    <= sub_wire11(3 DOWNTO 0);
	rx_syncstatus    <= sub_wire12(3 DOWNTO 0);
	tx_dataout    <= sub_wire13(3 DOWNTO 0);

	Hard_IP_x4_serdes_alt_c3gxb_41f8_component : Hard_IP_x4_serdes_alt_c3gxb_41f8
	GENERIC MAP (
		starting_channel_number => starting_channel_number
	)
	PORT MAP (
		cal_blk_clk => cal_blk_clk,
		fixedclk => fixedclk,
		gxb_powerdown => gxb_powerdown,
		pipe8b10binvpolarity => pipe8b10binvpolarity,
		pll_areset => pll_areset,
		pll_inclk => pll_inclk,
		powerdn => powerdn,
		reconfig_clk => reconfig_clk,
		reconfig_togxb => reconfig_togxb,
		rx_analogreset => rx_analogreset,
		rx_datain => rx_datain,
		rx_digitalreset => rx_digitalreset,
		rx_elecidleinfersel => rx_elecidleinfersel,
		tx_ctrlenable => tx_ctrlenable,
		tx_datain => tx_datain,
		tx_detectrxloop => tx_detectrxloop,
		tx_digitalreset => tx_digitalreset,
		tx_forcedispcompliance => tx_forcedispcompliance,
		tx_forceelecidle => tx_forceelecidle,
		coreclkout => sub_wire0,
		hip_tx_clkout => sub_wire1,
		pipedatavalid => sub_wire2,
		pipeelecidle => sub_wire3,
		pipephydonestatus => sub_wire4,
		pipestatus => sub_wire5,
		pll_locked => sub_wire6,
		reconfig_fromgxb => sub_wire7,
		rx_ctrldetect => sub_wire8,
		rx_dataout => sub_wire9,
		rx_freqlocked => sub_wire10,
		rx_patterndetect => sub_wire11,
		rx_syncstatus => sub_wire12,
		tx_dataout => sub_wire13
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: PRIVATE: IP_MODE STRING "PCIE_HIP_8"
-- Retrieval info: PRIVATE: LOCKDOWN_EXCL STRING "PCIE"
-- Retrieval info: PRIVATE: NUM_KEYS NUMERIC "0"
-- Retrieval info: PRIVATE: RECONFIG_PROTOCOL STRING "BASIC"
-- Retrieval info: PRIVATE: RECONFIG_SUBPROTOCOL STRING "none"
-- Retrieval info: PRIVATE: RX_ENABLE_DC_COUPLING STRING "false"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE STRING "2500"
-- Retrieval info: PRIVATE: WIZ_BASE_DATA_RATE_ENABLE STRING "0"
-- Retrieval info: PRIVATE: WIZ_DATA_RATE STRING "2500"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INCLK_FREQ_ARRAY STRING "100 100 100 100 100 100 100 100 100 100 100 100 100 100 100 100 100 100 100 100"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A STRING "2000"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_A_UNIT STRING "Mbps"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B STRING "100"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_B_UNIT STRING "MHz"
-- Retrieval info: PRIVATE: WIZ_DPRIO_INPUT_SELECTION NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_FREQ STRING "100.0"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK0_PROTOCOL STRING "PCI Express (PIPE)"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK1_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK2_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK3_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK4_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK5_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_FREQ STRING "250"
-- Retrieval info: PRIVATE: WIZ_DPRIO_REF_CLK6_PROTOCOL STRING "Basic"
-- Retrieval info: PRIVATE: WIZ_ENABLE_EQUALIZER_CTRL NUMERIC "1"
-- Retrieval info: PRIVATE: WIZ_EQUALIZER_CTRL_SETTING NUMERIC "1"
-- Retrieval info: PRIVATE: WIZ_FORCE_DEFAULT_SETTINGS NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_INCLK_FREQ STRING "100.0"
-- Retrieval info: PRIVATE: WIZ_INCLK_FREQ_ARRAY STRING "100.0 125.0"
-- Retrieval info: PRIVATE: WIZ_INPUT_A STRING "2500"
-- Retrieval info: PRIVATE: WIZ_INPUT_A_UNIT STRING "Mbps"
-- Retrieval info: PRIVATE: WIZ_INPUT_B STRING "100.0"
-- Retrieval info: PRIVATE: WIZ_INPUT_B_UNIT STRING "MHz"
-- Retrieval info: PRIVATE: WIZ_INPUT_SELECTION NUMERIC "0"
-- Retrieval info: PRIVATE: WIZ_PROTOCOL STRING "PCI Express (PIPE)"
-- Retrieval info: PRIVATE: WIZ_SUBPROTOCOL STRING "Gen 1-x4"
-- Retrieval info: PRIVATE: WIZ_WORD_ALIGN_FLIP_PATTERN STRING "0"
-- Retrieval info: PARAMETER: STARTING_CHANNEL_NUMBER NUMERIC "0"
-- Retrieval info: CONSTANT: EFFECTIVE_DATA_RATE STRING "2500 Mbps"
-- Retrieval info: CONSTANT: ENABLE_LC_TX_PLL STRING "false"
-- Retrieval info: CONSTANT: ENABLE_PLL_INCLK_ALT_DRIVE_RX_CRU STRING "true"
-- Retrieval info: CONSTANT: ENABLE_PLL_INCLK_DRIVE_RX_CRU STRING "true"
-- Retrieval info: CONSTANT: EQUALIZER_DCGAIN_SETTING NUMERIC "1"
-- Retrieval info: CONSTANT: GEN_RECONFIG_PLL STRING "false"
-- Retrieval info: CONSTANT: GX_CHANNEL_TYPE STRING ""
-- Retrieval info: CONSTANT: INPUT_CLOCK_FREQUENCY STRING "100.0 MHz"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV GX"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_SPEED_GRADE STRING "6"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_VARIANT STRING "ANY"
-- Retrieval info: CONSTANT: LOOPBACK_MODE STRING "none"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "alt_c3gxb"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "4"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "duplex"
-- Retrieval info: CONSTANT: PLL_BANDWIDTH_TYPE STRING "Auto"
-- Retrieval info: CONSTANT: PLL_CONTROL_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: PLL_INCLK_PERIOD NUMERIC "10000"
-- Retrieval info: CONSTANT: PLL_PFD_FB_MODE STRING "internal"
-- Retrieval info: CONSTANT: PREEMPHASIS_CTRL_1STPOSTTAP_SETTING NUMERIC "1"
-- Retrieval info: CONSTANT: PROTOCOL STRING "pcie"
-- Retrieval info: CONSTANT: RECEIVER_TERMINATION STRING "oct_100_ohms"
-- Retrieval info: CONSTANT: RECONFIG_DPRIO_MODE NUMERIC "0"
-- Retrieval info: CONSTANT: RX_8B_10B_MODE STRING "normal"
-- Retrieval info: CONSTANT: RX_ALIGN_PATTERN STRING "0101111100"
-- Retrieval info: CONSTANT: RX_ALIGN_PATTERN_LENGTH NUMERIC "10"
-- Retrieval info: CONSTANT: RX_ALLOW_ALIGN_POLARITY_INVERSION STRING "false"
-- Retrieval info: CONSTANT: RX_ALLOW_PIPE_POLARITY_INVERSION STRING "true"
-- Retrieval info: CONSTANT: RX_BITSLIP_ENABLE STRING "false"
-- Retrieval info: CONSTANT: RX_BYTE_ORDERING_MODE STRING "NONE"
-- Retrieval info: CONSTANT: RX_CHANNEL_BONDING STRING "x4"
-- Retrieval info: CONSTANT: RX_CHANNEL_WIDTH NUMERIC "8"
-- Retrieval info: CONSTANT: RX_COMMON_MODE STRING "0.82v"
-- Retrieval info: CONSTANT: RX_CRU_INCLOCK0_PERIOD NUMERIC "10000"
-- Retrieval info: CONSTANT: RX_DATAPATH_PROTOCOL STRING "pipe"
-- Retrieval info: CONSTANT: RX_DATA_RATE NUMERIC "2500"
-- Retrieval info: CONSTANT: RX_DATA_RATE_REMAINDER NUMERIC "0"
-- Retrieval info: CONSTANT: RX_DIGITALRESET_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: RX_ENABLE_BIT_REVERSAL STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_LOCK_TO_DATA_SIG STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_LOCK_TO_REFCLK_SIG STRING "false"
-- Retrieval info: CONSTANT: RX_ENABLE_SELF_TEST_MODE STRING "false"
-- Retrieval info: CONSTANT: RX_FORCE_SIGNAL_DETECT STRING "false"
-- Retrieval info: CONSTANT: RX_PPMSELECT NUMERIC "8"
-- Retrieval info: CONSTANT: RX_RATE_MATCH_FIFO_MODE STRING "normal"
-- Retrieval info: CONSTANT: RX_RATE_MATCH_PATTERN1 STRING "11010000111010000011"
-- Retrieval info: CONSTANT: RX_RATE_MATCH_PATTERN2 STRING "00101111000101111100"
-- Retrieval info: CONSTANT: RX_RATE_MATCH_PATTERN_SIZE NUMERIC "20"
-- Retrieval info: CONSTANT: RX_RUN_LENGTH NUMERIC "40"
-- Retrieval info: CONSTANT: RX_RUN_LENGTH_ENABLE STRING "true"
-- Retrieval info: CONSTANT: RX_SIGNAL_DETECT_THRESHOLD NUMERIC "4"
-- Retrieval info: CONSTANT: RX_USE_ALIGN_STATE_MACHINE STRING "true"
-- Retrieval info: CONSTANT: RX_USE_CLKOUT STRING "false"
-- Retrieval info: CONSTANT: RX_USE_CORECLK STRING "false"
-- Retrieval info: CONSTANT: RX_USE_DESERIALIZER_DOUBLE_DATA_MODE STRING "false"
-- Retrieval info: CONSTANT: RX_USE_DESKEW_FIFO STRING "false"
-- Retrieval info: CONSTANT: RX_USE_DOUBLE_DATA_MODE STRING "false"
-- Retrieval info: CONSTANT: RX_USE_PIPE8B10BINVPOLARITY STRING "true"
-- Retrieval info: CONSTANT: RX_USE_RATE_MATCH_PATTERN1_ONLY STRING "false"
-- Retrieval info: CONSTANT: TRANSMITTER_TERMINATION STRING "oct_100_ohms"
-- Retrieval info: CONSTANT: TX_8B_10B_MODE STRING "normal"
-- Retrieval info: CONSTANT: TX_ALLOW_POLARITY_INVERSION STRING "false"
-- Retrieval info: CONSTANT: TX_CHANNEL_BONDING STRING "x4"
-- Retrieval info: CONSTANT: TX_CHANNEL_WIDTH NUMERIC "8"
-- Retrieval info: CONSTANT: TX_CLKOUT_WIDTH NUMERIC "4"
-- Retrieval info: CONSTANT: TX_COMMON_MODE STRING "0.65v"
-- Retrieval info: CONSTANT: TX_DATA_RATE NUMERIC "2500"
-- Retrieval info: CONSTANT: TX_DATA_RATE_REMAINDER NUMERIC "0"
-- Retrieval info: CONSTANT: TX_DIGITALRESET_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: TX_ENABLE_BIT_REVERSAL STRING "false"
-- Retrieval info: CONSTANT: TX_ENABLE_SELF_TEST_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_PLL_BANDWIDTH_TYPE STRING "Auto"
-- Retrieval info: CONSTANT: TX_PLL_INCLK0_PERIOD NUMERIC "10000"
-- Retrieval info: CONSTANT: TX_PLL_TYPE STRING "CMU"
-- Retrieval info: CONSTANT: TX_SLEW_RATE STRING "low"
-- Retrieval info: CONSTANT: TX_TRANSMIT_PROTOCOL STRING "pipe"
-- Retrieval info: CONSTANT: TX_USE_CORECLK STRING "false"
-- Retrieval info: CONSTANT: TX_USE_DOUBLE_DATA_MODE STRING "false"
-- Retrieval info: CONSTANT: TX_USE_SERIALIZER_DOUBLE_DATA_MODE STRING "false"
-- Retrieval info: CONSTANT: USE_CALIBRATION_BLOCK STRING "true"
-- Retrieval info: CONSTANT: VOD_CTRL_SETTING NUMERIC "4"
-- Retrieval info: CONSTANT: coreclkout_control_width NUMERIC "1"
-- Retrieval info: CONSTANT: elec_idle_infer_enable STRING "false"
-- Retrieval info: CONSTANT: enable_0ppm STRING "false"
-- Retrieval info: CONSTANT: equalization_setting NUMERIC "5"
-- Retrieval info: CONSTANT: gxb_powerdown_width NUMERIC "1"
-- Retrieval info: CONSTANT: hip_enable STRING "true"
-- Retrieval info: CONSTANT: iqtxrxclk_allowed STRING ""
-- Retrieval info: CONSTANT: number_of_quads NUMERIC "1"
-- Retrieval info: CONSTANT: pll_divide_by STRING "2"
-- Retrieval info: CONSTANT: pll_multiply_by STRING "25"
-- Retrieval info: CONSTANT: reconfig_calibration STRING "true"
-- Retrieval info: CONSTANT: reconfig_fromgxb_port_width NUMERIC "5"
-- Retrieval info: CONSTANT: reconfig_pll_control_width NUMERIC "1"
-- Retrieval info: CONSTANT: reconfig_togxb_port_width NUMERIC "4"
-- Retrieval info: CONSTANT: rx_cdrctrl_enable STRING "true"
-- Retrieval info: CONSTANT: rx_deskew_pattern STRING "0"
-- Retrieval info: CONSTANT: rx_dwidth_factor NUMERIC "1"
-- Retrieval info: CONSTANT: rx_enable_second_order_loop STRING "false"
-- Retrieval info: CONSTANT: rx_loop_1_digital_filter NUMERIC "8"
-- Retrieval info: CONSTANT: rx_signal_detect_loss_threshold STRING "3"
-- Retrieval info: CONSTANT: rx_signal_detect_valid_threshold STRING "14"
-- Retrieval info: CONSTANT: rx_use_external_termination STRING "false"
-- Retrieval info: CONSTANT: rx_word_aligner_num_byte NUMERIC "1"
-- Retrieval info: CONSTANT: top_module_name STRING "Hard_IP_x4_serdes"
-- Retrieval info: CONSTANT: tx_bitslip_enable STRING "FALSE"
-- Retrieval info: CONSTANT: tx_dwidth_factor NUMERIC "1"
-- Retrieval info: CONSTANT: tx_use_external_termination STRING "false"
-- Retrieval info: USED_PORT: cal_blk_clk 0 0 0 0 INPUT NODEFVAL "cal_blk_clk"
-- Retrieval info: USED_PORT: coreclkout 0 0 1 0 OUTPUT NODEFVAL "coreclkout[0..0]"
-- Retrieval info: USED_PORT: fixedclk 0 0 0 0 INPUT NODEFVAL "fixedclk"
-- Retrieval info: USED_PORT: gxb_powerdown 0 0 1 0 INPUT NODEFVAL "gxb_powerdown[0..0]"
-- Retrieval info: USED_PORT: hip_tx_clkout 0 0 4 0 OUTPUT NODEFVAL "hip_tx_clkout[3..0]"
-- Retrieval info: USED_PORT: pipe8b10binvpolarity 0 0 4 0 INPUT NODEFVAL "pipe8b10binvpolarity[3..0]"
-- Retrieval info: USED_PORT: pipedatavalid 0 0 4 0 OUTPUT NODEFVAL "pipedatavalid[3..0]"
-- Retrieval info: USED_PORT: pipeelecidle 0 0 4 0 OUTPUT NODEFVAL "pipeelecidle[3..0]"
-- Retrieval info: USED_PORT: pipephydonestatus 0 0 4 0 OUTPUT NODEFVAL "pipephydonestatus[3..0]"
-- Retrieval info: USED_PORT: pipestatus 0 0 12 0 OUTPUT NODEFVAL "pipestatus[11..0]"
-- Retrieval info: USED_PORT: pll_areset 0 0 1 0 INPUT NODEFVAL "pll_areset[0..0]"
-- Retrieval info: USED_PORT: pll_inclk 0 0 1 0 INPUT NODEFVAL "pll_inclk[0..0]"
-- Retrieval info: USED_PORT: pll_locked 0 0 1 0 OUTPUT NODEFVAL "pll_locked[0..0]"
-- Retrieval info: USED_PORT: powerdn 0 0 8 0 INPUT NODEFVAL "powerdn[7..0]"
-- Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
-- Retrieval info: USED_PORT: reconfig_fromgxb 0 0 5 0 OUTPUT NODEFVAL "reconfig_fromgxb[4..0]"
-- Retrieval info: USED_PORT: reconfig_togxb 0 0 4 0 INPUT NODEFVAL "reconfig_togxb[3..0]"
-- Retrieval info: USED_PORT: rx_analogreset 0 0 1 0 INPUT NODEFVAL "rx_analogreset[0..0]"
-- Retrieval info: USED_PORT: rx_ctrldetect 0 0 4 0 OUTPUT NODEFVAL "rx_ctrldetect[3..0]"
-- Retrieval info: USED_PORT: rx_datain 0 0 4 0 INPUT NODEFVAL "rx_datain[3..0]"
-- Retrieval info: USED_PORT: rx_dataout 0 0 32 0 OUTPUT NODEFVAL "rx_dataout[31..0]"
-- Retrieval info: USED_PORT: rx_digitalreset 0 0 1 0 INPUT NODEFVAL "rx_digitalreset[0..0]"
-- Retrieval info: USED_PORT: rx_elecidleinfersel 0 0 12 0 INPUT NODEFVAL "rx_elecidleinfersel[11..0]"
-- Retrieval info: USED_PORT: rx_freqlocked 0 0 4 0 OUTPUT NODEFVAL "rx_freqlocked[3..0]"
-- Retrieval info: USED_PORT: rx_patterndetect 0 0 4 0 OUTPUT NODEFVAL "rx_patterndetect[3..0]"
-- Retrieval info: USED_PORT: rx_syncstatus 0 0 4 0 OUTPUT NODEFVAL "rx_syncstatus[3..0]"
-- Retrieval info: USED_PORT: tx_ctrlenable 0 0 4 0 INPUT NODEFVAL "tx_ctrlenable[3..0]"
-- Retrieval info: USED_PORT: tx_datain 0 0 32 0 INPUT NODEFVAL "tx_datain[31..0]"
-- Retrieval info: USED_PORT: tx_dataout 0 0 4 0 OUTPUT NODEFVAL "tx_dataout[3..0]"
-- Retrieval info: USED_PORT: tx_detectrxloop 0 0 4 0 INPUT NODEFVAL "tx_detectrxloop[3..0]"
-- Retrieval info: USED_PORT: tx_digitalreset 0 0 1 0 INPUT NODEFVAL "tx_digitalreset[0..0]"
-- Retrieval info: USED_PORT: tx_forcedispcompliance 0 0 4 0 INPUT NODEFVAL "tx_forcedispcompliance[3..0]"
-- Retrieval info: USED_PORT: tx_forceelecidle 0 0 4 0 INPUT NODEFVAL "tx_forceelecidle[3..0]"
-- Retrieval info: CONNECT: @cal_blk_clk 0 0 0 0 cal_blk_clk 0 0 0 0
-- Retrieval info: CONNECT: @fixedclk 0 0 0 0 fixedclk 0 0 0 0
-- Retrieval info: CONNECT: @gxb_powerdown 0 0 1 0 gxb_powerdown 0 0 1 0
-- Retrieval info: CONNECT: @pipe8b10binvpolarity 0 0 4 0 pipe8b10binvpolarity 0 0 4 0
-- Retrieval info: CONNECT: @pll_areset 0 0 1 0 pll_areset 0 0 1 0
-- Retrieval info: CONNECT: @pll_inclk 0 0 1 0 pll_inclk 0 0 1 0
-- Retrieval info: CONNECT: @powerdn 0 0 8 0 powerdn 0 0 8 0
-- Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
-- Retrieval info: CONNECT: @reconfig_togxb 0 0 4 0 reconfig_togxb 0 0 4 0
-- Retrieval info: CONNECT: @rx_analogreset 0 0 1 0 rx_analogreset 0 0 1 0
-- Retrieval info: CONNECT: @rx_datain 0 0 4 0 rx_datain 0 0 4 0
-- Retrieval info: CONNECT: @rx_digitalreset 0 0 1 0 rx_digitalreset 0 0 1 0
-- Retrieval info: CONNECT: @rx_elecidleinfersel 0 0 12 0 rx_elecidleinfersel 0 0 12 0
-- Retrieval info: CONNECT: @tx_ctrlenable 0 0 4 0 tx_ctrlenable 0 0 4 0
-- Retrieval info: CONNECT: @tx_datain 0 0 32 0 tx_datain 0 0 32 0
-- Retrieval info: CONNECT: @tx_detectrxloop 0 0 4 0 tx_detectrxloop 0 0 4 0
-- Retrieval info: CONNECT: @tx_digitalreset 0 0 1 0 tx_digitalreset 0 0 1 0
-- Retrieval info: CONNECT: @tx_forcedispcompliance 0 0 4 0 tx_forcedispcompliance 0 0 4 0
-- Retrieval info: CONNECT: @tx_forceelecidle 0 0 4 0 tx_forceelecidle 0 0 4 0
-- Retrieval info: CONNECT: coreclkout 0 0 1 0 @coreclkout 0 0 1 0
-- Retrieval info: CONNECT: hip_tx_clkout 0 0 4 0 @hip_tx_clkout 0 0 4 0
-- Retrieval info: CONNECT: pipedatavalid 0 0 4 0 @pipedatavalid 0 0 4 0
-- Retrieval info: CONNECT: pipeelecidle 0 0 4 0 @pipeelecidle 0 0 4 0
-- Retrieval info: CONNECT: pipephydonestatus 0 0 4 0 @pipephydonestatus 0 0 4 0
-- Retrieval info: CONNECT: pipestatus 0 0 12 0 @pipestatus 0 0 12 0
-- Retrieval info: CONNECT: pll_locked 0 0 1 0 @pll_locked 0 0 1 0
-- Retrieval info: CONNECT: reconfig_fromgxb 0 0 5 0 @reconfig_fromgxb 0 0 5 0
-- Retrieval info: CONNECT: rx_ctrldetect 0 0 4 0 @rx_ctrldetect 0 0 4 0
-- Retrieval info: CONNECT: rx_dataout 0 0 32 0 @rx_dataout 0 0 32 0
-- Retrieval info: CONNECT: rx_freqlocked 0 0 4 0 @rx_freqlocked 0 0 4 0
-- Retrieval info: CONNECT: rx_patterndetect 0 0 4 0 @rx_patterndetect 0 0 4 0
-- Retrieval info: CONNECT: rx_syncstatus 0 0 4 0 @rx_syncstatus 0 0 4 0
-- Retrieval info: CONNECT: tx_dataout 0 0 4 0 @tx_dataout 0 0 4 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL Hard_IP_x4_serdes.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Hard_IP_x4_serdes.ppf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Hard_IP_x4_serdes.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Hard_IP_x4_serdes.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Hard_IP_x4_serdes.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Hard_IP_x4_serdes_inst.vhd FALSE
